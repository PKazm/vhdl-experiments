// ********************************************************************/ 
// Microsemi Corporation Proprietary and Confidential 
// Copyright 2018 Microsemi Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
// ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE APPROVED 
// IN ADVANCE IN WRITING.  
//  
// Description:  Block computes:
//                 1. Natural log of a number
//                 2. Square root of a number
//                 The block instantiates a hyperbolic CORDIC block, and 
//                 scales the result appropriately. The CORDIC architecture can
//                 be selected as:
//                 G_ARCHITECTURE = 0 --> Sequential
//                 G_ARCHITECTURE = 1 --> Pipeline  
//
// Revision Information:
// Date     Description
// 07Mar18 Initial Release 
//
// SVN Revision Information:
// SVN $Revision: $
// SVN $Date: $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes: 
//        
// *********************************************************************/ 

//=================================================================================================
// CoreLNSQRT module declaration
//=================================================================================================
module CORELNSQRT
#(
// Generic list
    // Specifies the type of architecture(Sequential = 0, Pipeline = 1).
	parameter G_ARCHITECTURE                  = 0,
	
	// Specifies the input bit width.
	parameter G_INPUT_WIDTH                   = 18,
	
	// Specifies the output bit width.
	parameter G_OUTPUT_WIDTH                  = 64,
	
	// Specifies the number of iterations.
	parameter G_NO_OF_ITERATIONS              = 25
)
 (
// Port list
    // System reset
	input RESETN_I,

    // System clock
	input SYS_CLK_I,

    // Start signal for cordic operation
	input START_I,

    // Input
	input  [G_INPUT_WIDTH-1:0] INPUT_I,

    // Signal specifies cordic has finished its operation
    output wire DONE_O,

    // Natural log output
    output wire [G_OUTPUT_WIDTH-1:0] LOG_O,

    // Square root output
	output wire [G_OUTPUT_WIDTH-1:0] SQ_ROOT_O
);


//=================================================================================================
// Synthesis Attributes
//=================================================================================================
//NA//
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="author-a", author_info="author-a-details"
`pragma protect encrypt_agent="encryptP1735.pl", encrypt_agent_info="Synplify encryption scripts"

`pragma protect key_keyowner="Synplicity", key_keyname="SYNP05_001", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_block
e+LgDzWtd0Y6z2rbdVcAuFIhrtPrbjoDvW2SFEvNPAF2CNm7QvSVaYy8iqSCVI3DSqmgPMjc1Vps
8uvEH50D1YTwO0l0Pw75Plb8lhq8MsMg7Z5FzgynoBRft2eS1C/KpF2ixqe+Zo9ynavI5TR1wBGo
MhkfjqNMAh5e8eVLHoAQ9XL/OND7Jq1BoL+70hz+8VJSoxkFhObF9CV4qrnpJJt/VI2R+Slzpd1W
oFtfvvkaeObq8tIpYV6eeNMqsS3SGx+x9GExOh/mVeUIqi9hWmVizvDUs12X04Ube8bYNlHfNIJ4
VqWuPdWAsGC/+lw1XaH4EzjZyaXLncPpwEKWEQ==

`pragma protect key_keyowner="Mentor Graphics Corporation", key_keyname="MGC-VERIF-SIM-RSA-1", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=128)
`pragma protect key_block
cy+Big5bidjybxB3hnsXKDaHMHwYklHNuGf6tzhD/E3Bz5AkbzJYcq6nXNJXS7MR9vA56dJ/6vB9
EXkAlGQvgtx519NuyFFiG7cgN48rGTGbW5COTub4Jk2GeD+IDviaCPoUNMxDfu/g64zwAA0Z5Vyh
UaiWxEhb/xw0h3/LFOA=

`pragma protect key_keyowner="Microsemi Corporation", key_keyname="MSC-IP-KEY-RSA", key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=960)
`pragma protect key_block
N3/aD0M40ObkNHQ2rCtrgYgPNrrH79UqhrY+JIRCSAaLo19QbHpzGuu8EktpnxPw0kELwEpL8mjz
aeob59EGxGpJMk8OC6FBvt0JG8OWVlqAtYlidpuO6CfO3TW+okLzNwjD+1JrTu686lOjfhTfdsdJ
8qOS1ZNat9gPwFabYn4Xjs8x0G/2w9ku54+2tXDuSG3LagSQtuUWQCwhj3oZnypaB0NpRfc1rn+W
6C1+q/1iPh6IiGSKjHkTASKXknlp7xVFnGNe+pNR192QUjzWDHWaEhG5hGWFo5NaCX+zFkbJHe6C
b7aZVssdsAEHivZpifM+bNt8PGI5+fYFnNpgN+uGgrA3e9OvcpHfpgKZ6XPjGSgvTIBNajSGtvtD
ynaNXESL9HYTmOHXdSUerrwXLNHzjNnrJMpVZBv6zKlkVt1K8XmNxOnssVvTQUjdTMNVmZvwuhDo
vAn27AEmIcMq5mZeGVA1agRoG3IrL0KQWk3RJEzt24G/PCBiB70Sl7DTG6/e6hBeRUPOG3oIG1Cq
dMcOGr4QVXogQl0Dql9ubGqIzSU1nGDuwgMwH7SpB9utkGYBkaxNQZpagnLKi9srTDILqdd1GuYC
P7VotT4o2FcRAvQAvRVF80iaW4AdaoMvnbI4+p1qwsN+qd800iEBmPBUSZlHQ1mKuGU758rczzOI
zk9/ZGeCFEgApKeCiD+8IaUjOeNtCGIJ55VNQFRZtAUbOR1X9DKuXRM7wPYQvZCqQDI9zOweEvoI
e1nnE5oWpwg69kd2CoDMV9n5fX39NXaOQTqE/nrOkib2gQbev9quCVz84sSSy5HXp8XrFs2C3XDv
aaXhHU+rX2Tnc/DadAc72pYkR2JXUWUUrdcHZCvl1Yv5hMW1lx/mbRM2CAZ9jLrP8lfT/DzXWFX2
kU+5s1BbTDlKOtW5w+USS/5DOwfjeS76ifNAWa/ffsi77hWi2rf8rTRCQteulPulyDQf5nULP1GV
drkjP5K6wq2suau2a+igPT9/khD2nxoNM0cEhZsxIyUp1LUR7PdFRm08gCuuijWcpXEBUQHwWwbk
zFqhy0JrA9MGSLF0UWrwb2JAZATg4aTZmwscmRbU5rZozSI3Wa+yBdt5QRQhfCdOuiOc8XZQ93Tl
YAOJ9nOb5CedAW9Hy+iEtOBem2/Xha0L5q8QOBjV3L5PJY1yO7qr41jkuGSZYnNl40ccvI2WYYul
mKDU9JYMcv0qv2bkYpzBFagDkKEC54J/U17/7X/rKpzb/nvA/WZWPrI6HaIz4lLX

`pragma protect data_keyowner="ip-vendor-a", data_keyname="fpga-ip", data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=44896)
`pragma protect data_block
a4DYV7ZfIiHeTXYbab9UGzTnE3RpxKC5aGOCXOpofoN2pL9orY1+iBApnvo71L79zTEUw5ZfAjEo
GXAb8ZY15Yt8BlYfPek9tH2i7zYKc9VtrH9Z0KIvC9rnZxG0ha3/XGQKsu8zrR6PMXgSTlgrVq6j
jl5F/JrKrdu/1Vg/mpX6kniTGpd67UhBM5sQ/6hz7T/q72aAFI76xqQOgRLpdABzH5T1EYEH+ifi
UqPcrT3soi46nwL9HhkKXVjPRGLPfWro8hVF9ywjeVH/pJW+YwUs8NOOqXpyybLMo/hBal+Wx5Pf
6dVyVJOwYbNe3q2uXUd0+GuZZX/9jR93GP6FuqXivnffDZooBURQygC5456ndGruZOW5bBt4he/P
U48dqzel9O+pT47neMVW0mJqGXPgB9idgntTM/c3fgIZPmstBzuesfkdd+ikuij7N5MFDWIehZYP
ERHK0R1k2KJmVTFqQNi+BepwN+J9F3+g8Y06J6HZxjbBan2gq6DBYvsxHqcURl86XfVPdber+AQ/
osJilD32H2IDkj5yLQ1OltLA0qZqSC3phk0MV5kyC4Z0ZSHyIKks7VjqD3hZ9Uouaj18rZP+lxHB
sV2nQq329GuetDSgTmHKbj59IT5hKbe0/5/GYcMNnv86vDuwHH18BUGrkeGd4EDXPs9gK0AtWeuq
ovN7fr2DhCZaFXdEDx8tCCkcQ1qknSKVlJlZF8ZhGDPgQYisrNTRXwExxzhSh6Kufl39jhehXPHz
yIRA96U7lvCcoDUcgqvSeZQ4ucLyJgV2vob4VYJzOKwYfP2dCIBgtBbsCOQnFytPluCHSHDyrvlz
lPH/hLotfPjhT42tsFUoqQPnso5XdXoBxuFQh/DR0qZE91yqjm9d9lod26cLdoGpER8ulZICbE1Y
3RvJjGg5jjwlW3KrdgHCC+++4ycc/LaactyZYGXdcMUjIg2+qrgqNrWdYmHC0DiVlRw3nq/yXY1v
kTsBUv5X8LBb0nTuN4kgoLtRkSi7XQ3eJeUMECASgRu4ntCZ1PpSgPqm+7Psni1dCBDe5YoWjwCQ
BRJ88JiGLgnfThjJzUfVvdwrdQYQ/us91dgvTK3iNGFE6YuO6rs22eWavvlzU7Yko2v+HltUSBHc
gmUa+dq1fG4v5p15IomMGiFIQTy5CH1qqcC9ZfTxXCM1aefvEzQ6I3nUPrHruC3c4N5YO1ztIRyV
9XBrB8NGmdPr6cIPU1gkhKFdI08Ovf8SryRoyeDl6Lk2w7WBYgk1qjC+n2iCkvh4zjy6v5bJKhvB
aXlr2vxCDdV9O3r/5fSqyxQ9QwZS3FHevgIbrLmlXgHjZJtoz4DtO2FenVpOqqOCLueiir73jh0q
SkEps+tK36QylOeSc2IBFzY6Bl8vEXXTkUtLrpbPmlGdf4WYlKOcJlE0QwDRac2VSHfG7d/B6bHI
u3Mga/e83F3O15L2INSRGXNTCQOPywcNnyf4q6fD7LJK/1Sov5ix5MRLMhArDyowgQNB1hoiKpv7
CBX+fdZW8F3yaNyPRjzeaRT1qg9hOUOC3QKNnuG2WrGflZql3wGjvmkn4MQ0P3JKwzHpI3MBvJH9
MuT/QVq7SOJ6/yG4On7vLWlpZHiCxQN03FtcIUYEKoXy9pG7RVv4SRpiUbMFkO7YnVGFx8pNCfHP
3wSUwvhzXJB38ynFfE/CIzLXpJgyuOSYeInHCJkZHEoOpkurpQXrJ7zrWmQXX3FHHI2te9TDJJJy
OJi5HJn15J0H80MYpyOLIHEzZl7zcKQk5oFxn6YjIW0UMDi+YfI3vJ1zks5GRNPJBGD/0dA15oJD
pT488dRxN/+CxPkpVkvWV55uOAvJA+WC72ybSi/Kv6ughEHirmqdD6oime4qutcuM0KnvCzroIZD
OAY01wXF3TGolhk1Utd3Disaa9ElCpVdMiJ7LL35y7rKhZVPYgjl3mHgHYFGIGKmQIvstrGAqTe/
iWJ73jHp+pKSnyUPSX2XrnUdMMJP/OnKYfiKA23jNpVfiGhOZBCXLXBLokG8XyyX7XMY65q6TmZS
kGax6djAKwsl17DAPYXPZnkl4/ACBjizHo/nmCovERqMfXBUK3lFqhsDo15Q1yyZ+C5u5/v1Tdj7
X9rUaO6aK1w/N3Z10xxGFK0vNxusOd9rnYC8CDLBwgjvFSC+rhZTc1OTSXuhlb0UMUn0YaebKcgU
yVnwDx/Gow+3CPdwSX658D61MpOou5s9pblQvrfPYqVt562pCWWU5Nh4kRV4Ym2zAlr8WPeOZ+fQ
vamJ4ep4QuGCHB+PyGh+tpnoA62hmXyL+wPGpdIC+8kY9Xos+yU+D3zRl1Vl9tsjEwS4pauWXZny
Yi6hr5UYHodHgimiC9P/vI0iNjiqi3JG1mdkZY82H0ohLqwIii5o+nJbhDDg4YH5V5+PjQgZ1iQo
Lj9scfvBmP61fEu4ea61zLes6DbBGuQtpLgZHE4nzDd80QoaiTpt9MGegn64+vTkUeXqLx1Z+n/R
dyLIWM5OT/WVUglRNHlPvwPxSPGXdN0582/Vv+Ntmsbh4yz8qMO11k4Tpava1EHJd2LXQs4+0+sw
Y4+lBq+JBc2vrWGKU1ChqsrdVwvbeNkqBTa+KIcQKcihDeZ6YhHh4pR7wZCl6bTMxpHv8BcDjRZU
sDhYFtOxNeBnwQyGBMt608Tjdnd6bh1oo+r8zTV5yHc2BAOoEO9bY1fFexWdcUpQUuIu7x7fnDso
dJ4GHUZzMxObIZCPYDWc9YrEM+OHeVfmVNvhYX4Hr17GNLZoacIndI4WwOA4C7bsUVfkYLTyRewC
GgAo59zvrRJTzNTeBnrlwbO8RMi5S1i9LgqeZmiBsDf1wkNitlHPb6OqVL+7U3zDQhQrkSm7EGKC
wqlXCjWFAMxlyrMYYsbi7H8JXK/TP+UgYJjLHFI6bdsGTmW000nOL31HnBBmJMW0rlq1kfGWZtsc
lHzqVti61AMpDBc6GSKs1ZYALSed6mgm9BBgDVsw1y4TA9OlADpciBKJuKpwlD/QsA9hE0P558Xa
5BvWdd0aEVuktmiwQByDURAb9X+dKnCwCoYlFZkXT/zUW+Cm4WWBGOObG+llxAvNEXIob2TTWGMw
Ta4UKAIbKNOoUaslhARnBV9mFJc/hKosB8r6352XVvEePlBkhdnasW9RaAPwm8sLim+EBx0cfswi
woru+kF9/J5zdgQSdHFnHEO3R3TG4GEYko/TSKfvQn7Bck4E95hXW+12XOic83hAzVzleptVQF+T
H7Na86gW51tts+mNlmIZh58LI/273xGxs35ZOw6RmF+RyjrZ+5TbCrY7c02RQkcLCPhtUX/IibbD
xFJ6SpPzYVn+bhTGiwDJMbqciesDbhRl+nPS4Qkl0ugiPZyXqXguYgYMW7wg1dtjf8rl02PgMJLF
vg8EpIGN07KLcz+2N1F+xwvxvdYKj3x3gow0MsdvJ8OQ00vMRNkv5y7ZNdgLex2vLpMjGEgRZ495
0/ylvZT/WYCOEUWx/xwg5thBffHGt3zEPpG7p1s4AOApyvDbpLLfX6lkDAIkrBoULk1+EcP1ri5p
XbYvXzdw+TJvZi/10tIulE/4q6X4gu1f6PKYPp4TAlp3NaiVS3cnA+tMuiPE+J9+9kp51Tc9jNmz
iRz61T/KZewOfgdicn8huWaOuswtObxcfwsk6SMM/tzn7PDfN7IFsma7TBgGGkOaEs0A9MLSdBCs
cr/htw9NoCcJBbuiIsaXcxJcXRWZ+1FFqkd4gQWZGjZd/oYrQrKeY4aPu5+O0Y7HwusoDPwYMxxz
5cIvST9dvDcz1TVivpYqc9g4nYFBeWhD1M9tBURAEMgd4Ebbn7h3/P9T1nT9u5Xkws86ysbYAKGW
ygEeo7oaihJdG7dHISkmDr/mwCRxqiULTFklP+/LREWz1sXAgOzMgf2M6VTT46uy+13secdP8ImD
XBUg88XB0UVqU9ZyDiWun2R7biWrgeP1WVYgZ4OQmJtHFvvzEMcJEw7+h1AwqvCpSzPxj0M+K9eq
5Pj4Qvc8sqz7fkePhCvGX7I6bm9vZAjQ4savCxrWN5RdVbZ45r7EeGkOTle6NxvPoLQ2yVCUmT4h
v11Gflt52OHtkMa12b61IwwSQkZ0WzgXZalgdsLnva7TB78/T+yTvkvSIyvSOp7JFVq0BZyXaMeK
wyLE1z/BarFuyfuATaHAW8rH0Dhl6UHTVdZL+WcAA5SjQQxTtDC0nfMTKgtkJ/8tfwVyvbI1C8Fh
X/SpDHHnX7lKfn3F3lKdzrLSLxcy4NAOXf4OS6SalH0b1Db8AssmyMmVS9EYlxFP2q9lPCK/pLbv
1L6SJr3ipYnLfgkcDvVyOY5dIqWu4Cewf7q4i07C7HjXY4pxO41YCmBS4q5pmM8q3rCl1pl2FFIw
9/KzWCb+7q36QUTDTe92hOs1DqEcYIKnRYWZoBD3h5QLn6VPFbjeQwNwistv+oDhCd8xFJT76XO6
hB1zOLT7J4cHzCd5hn2MT6GCaPrqaOeNeXRs9Zqr22M1IhbzRV/fBYsNzD0aV87kumx8pVBo+wiT
L0iSwhGKK/AhBYDccE2M2gde/x47N7r83L4uqm3YcVG8ijvv/nCqCZo9T+sI5VKQRC3IzEw+MXTn
FoMUhwCrA4KFI3IVxb907rfdIThg5vSakTg7Eh7VuQP+ZmHrgO17dS6LQnplbM1nyTadDKHFjsF9
eI70mTuYOrXUXJPH9HjNjIgpz1lj/Av6BhAP8YO8oZD45y3J523NVk7o+ZWlEh0JVi4gRF9FQ8CY
rXPUqI0W1tHGQi6Im4sWRNVlz+qQFHIoRI2Zj5XWC41ooe074qj5HZptQJ9rRqj3T+KBlehGiyi9
30jGPFer+frK5NXLzRzW6s+u1W1Lz95ZHWW2kiotlmbTap/58FYRuDG4U2UIsnV07+JvUVTE+UmK
I/Pkbcl5YcoScmr5ESwLc5NNl9BAR0la1IvgoarMy0ImHesa59iE1BdaYUipWtUZlxwLO1yjmWgW
tGp7xP1rDbV6bA/3vRPdihOjlnOsMKcdM+/ltkvrZjC7EOp4/JqY5zVjMve3nigOu5k3kfyHJinr
ts3KkBepaN0Ld1ylR/G71Ipieft7qhFyXHv9WmH5fOby68/iJbgtypyXfLfvK0iW4rnqjUxGQTi2
kMy2MaUOQ7myuDitx2709kj6LDUUqHeQ9amArE6PxU+2XuEB46nL1T7c3vitL+3I/96AAyxjys9T
Mijw3L1ah0+U8RNoUIxj5cOSjSOCRdHaieEOc627fJCWuEQneDIXNj8OVVWaGRZQYL4aqcDVHq3b
XsDqtZ/hHuR6LLD1XKgftDyBCeeOA1/lzadwf7Sib2ix99ZDz3nfH1bQ1EWu5zqpADEEzec1OHwv
YV1AMiDM0cyrQZ97ul2G7654/RDY7rmgnxBGLbeX4d6TRUWbCaxLECd6Pj5m40i1xZl5hztnPFsC
tky/TJfXgDvVv3Eww5OjFvXlofDUSojGmll+qsDiH3NLwM+CJVHArKn82tAgfMTkHKXSfsavL60B
sC0wZt1tVsByoq5HnFGoZKrr/+6ura0cAniSyJQkoEXiqexN1WSiU4kkOUQpFZyOpErBSLY1/EBZ
+746zwQE+m71alEN3I/utFwlYD1INXdYexnTUUI0hLkjwljWuYOFx8Oxy450o9hhtuttPL1ILuAR
tvS5wTzrbeFuCNArgYieNNAFWTr0NgsGTi/S/PNTm4XSs70/dEP3mLWcU766K9UxRVxlgOcPibl0
N93GA25jwgDJhVO3skDx6E0bQWlZFE9tsPvdBdEBQU/zAM/kT4S9MfK9TdOQjuvi0U4pM32Irdzl
LnDUw4lTiaHp6wqds6WdunZmxqnyYXyDL1cq/S1gtpY8oyyTjzi9TOjso2UYgU9ryVOTeL0bY0v6
90VMCGWUvHBXkHZh5Zs+NIfo6k5dkXXyG/jWdDTVphBuxEB+2BUGfmrzG0dpCJoMAzBCqEb2IOK6
dhGWqfEIuFXo/xw4fKneuvkktPbCGKYN1CzddjA7gq2/zomJ6bT1ig5OT2vo88F/X0YNHNYDoc+P
M2sVwGfwsc98kLdolar1lJ0OWq5yhKDloR+v66jirtEvqvcGGXhNCkKVXWhRsc+8ORoV5iCUWGHk
QJWKAWDuJFbKB5+4WciuOyAf0m++iyn1EdLeXpEv/4C3CCmABWGq/JK5wKtCOHiTmVgKIOssD0sF
9KB1HdNbmPNy/PzAoE5J7qNDmzGgyBfHlfPz4CZklFLE3hSZPtXh+FnlnWA6AgMeelJwsCGYXmZi
Pyvj+Z0SJnlea/SlVweQ+k6JUoil9TtopNUMJisq5f0GW/2oR09xWPCp7rwP4qFSCAeFDOB87jNR
3F0KAwNoHYeyqr3KW1q8NA0JE+aX6mIHLRPZ0yl2Kts5VZro8kcLYezd/4k1SO3gobzq47cmJoTM
oUd8afnFIcpmGQ0dkEtPEZCXyQZksPxw1RO4QBNlwjGLZn8W1LpWkIj73B+BVSXCpW3YAHoTlY1M
M9BLpMOUxznl8Z6/40Y7jkapMxr3sbzueUsUzXSoM1DlTwdBN2VigvEtpEmipVTuXY7sA1+wS/gI
kDWLgHHfHONKLLlxsokpV8wL/H79Feu6sgm1ze2GL4+8wwHn77vwo2CjbceS1DGadkWut6xBI58D
nZRjwRZ04Gc1jzgubgS9WEMh17Fi/bhhn1iDXG1JwxecTJidKmDP5orbn0pDsg/4NqEZS5crPuZt
qyvJFZOOGABQPW4E8Z8axZ/NJi3IteW0wEzBuQR3r+8mVcBMgPhxlVvfvQVsLbLJ8mBTCvaAdA1e
kBSW4KRp3i6mSZ1QbGkMOId1DmZEgSChtPeFgNJf9QGqjFSSBCC5251FnDwf26ETuGsP4krAFDe2
VlqQidyTNk1tUtvyTMUsp+L6gIzEUrpDaBhpNlqSVHU+Fn5ziGQw3/hxNcNRtKvoUXHQQjTteWmT
CtrrLC/HxAYxHnywulI/6VoSlSrYo/AAp5UnKVjxu0gMB3yVG2eL8wHCyXB4000xwRoyWd8jVZsO
/fOVbzhyibjepMM9soHrMzahEhbEV7Tcgjhiyh0wCTJgmVOS4pwiyILziElSfgzeTTBrcloB8Gas
X3UTuG9JhXKruBOQ+Tt+UTUqvmxgJM+whFbK3vQ6a/TY4TCfy9uEJ1Jfyt9UVDtJaa8H0gx5Rmn0
ClIa2RdG/j4vjo0y8yHcBeL/y12EPBXpGtzrC/73GJYVpYlyxvL4bP8K4ae614XNEsT8ew0l8hRk
qPjdErcJmiJ2OQadMwqiCSbUTrYbIt/T3PfdDxBtMNzVRdO7tc1ZBWEnvZ+VOfT6/3Byl2jAfeON
loWXQVpMnsHm5BcPDBWckgstDo8JRmO7maFrHJj1MKKYNv91slQAoQDP89BRd9NO98TyNQ8dApD+
gIbo29zMa69oNKJVe+6f3wakP1P8eH//3PAmhZIPGUjmxJBjfFAq+/uzLWQTWbx26zNjUmNx9ziq
GIBofeYd/uE0wSw5hfqqMojbP6l8mT/2xqsYjVCZ5+cUNuM0NvR0/j14vWK/7swL/aH1Lw9Q+9e7
xPqjUIFXSSJG5WU14ygk8XxvCyRDItPfn5HyhCS6kyhhEBWdnsEGACRi7FuDvJPbtjO4ECJJ4wY7
DbEucjL2d7iKxG3HN/+5nlfgXsi9vsXnUWNZkzKdwglXuFWsXOHhENCYpzUl+ZN59AErST+fwpOH
3rxz9yWhDbj8QdujWR+Pos0eEDVVytPck8WTjM37QUqZANwR3+7CAdWvM5xThThXd76fJhVQaZsI
Q7EUbeU7lEgotwikW+DdORW9iFwlzlxBjKZ+Ejg+IeLj96xIq9MAnyiEoCeVRHHBqNaKyoAsepOc
rbANCU0FUrDi8g3ODUWi1wyOhDQgZNzhqRdw5AoXL+rkWptzubnsFI8AW8jWnyyKQgS0BgDpr7za
DWZ0WWIu4zs15KYAQQPHQZSE9IfBjnpgaz8xHuu7M1zcZGFKqSQUscG5Tr18H7gYx8In9XI2uEXk
iiwWngSOq5NdRhpTD4iJZq+TJr4TSE4Ztc099iEBd1J8IPouXGco1OcRkt0z7wGetuKTIJsDvq15
9ixkSvQXEUnPDO1IKWSQNW4S0WOk5XFhQKO64WrKbIdqKK/FXi42mqqL4pNQTvnyDL8DZJdbzwN+
45mOWieeXeWzvi//kIJIe4fWa7mKcBk32exga0/xZHVv/8u3b9iHg77Vc58iozr9Q3RhK5oAH2UI
IwLPugRHc6EUaP2xCaSVINVJzTSUAafJ88rCjDwT0Pr+QdLGfwGCBYPfknUYoQNM6jViK9WrBhU2
fNW2BmK5206jcmOF1qDrRfaGGhGkSkmnOQvgUslZDM74Dox7nyPD4NqMBMzGfmUphKeauOhIAk83
oavskyichhroIXxdWmb/kxNobY4kKOuIp0cKQoRDry99Ex9WCbFdC9tQ15PKJnzT37XuKLDBTmVQ
4zat+9p9P1CHWaDq6rqTBjgaBD3r9J/kPy6OvXkJQn4DdRncuVLtPBx3/+ubQK7EIAQ2f4adTH8Z
5KkGgC4Vu6HKQUahM1B9onvIj0j+VS3SUrRok3xaFPnh/ifDR+3NI0la+fi/tXpq0w5b2dzKQEEL
WXWt72mgFk1hoNaHRT/WYIKVfxPYmQItSzp3G3vRdRaDFhZqP167Ji/+9U3cEoV9ueemIT86UI9n
4mOWCjy540ZVifBhntmgzlo4svoV4TRDfeaeU+ihQJduz/LMM1ljf0KQYl2HkbNZlWEH08o5qi/G
7eznV+lrXhLHWhd//+ZK89h4I2OO95riW43V3Nu5xov6jHP2E2dZLJsnpIevdZKuGbVk9CZbsEZT
Nsd/KjMsLU6NIO/Xn9WGlj368PdLjZ6YCpWrETdB4mCjui2tK4h9aiu5pucqC0sVDiOZOWuHclNZ
/c4b8IJF2HHMZiZw8XJYLFCvy2939ag1uqOP583Tso5tSU9b5/UGkb6hCysXQkp/ssim57OH0VMO
htATK/LVReo/nSmxy9sU5DVn3+SepClMLVF9Q7UOcz1dZkkSpF2X8UQTfqWooFp8OKjPL9hHjehH
gFkb+YJDQ9xwB3Z3kXq2ztp37qDs6UEs//OmwOoAOvPOcFboIYFF6L283/oCArGQwwEgybOQQ/UD
auxIA7ri2UUXZV0jwlbMkBUXI0tNwSESWl/on20HqIb0mLbq8xLwJ2U9pkbp5u40gh+F8xp5H2+P
rHFo4Jgtnenu9cRch9F8kUJg8q2s6no+rJ6A4lFxUvnFI8/tsohbnDnXiSySZ23q3OC/+H1PD/sV
23ac7vRNbyHyedDy+4Sj6OAoNqAxPjZJ9g/5ZyzaDNNvsGMG93DTrCAzV4+iJha6/ksHOq9boxFu
rxwuGlaj4hpqKZNvwYSfMb9dIlZuMhvXMxS+mZ8BLEAT5gFCyPpmJYYnQf69BHyT8gB71yz4ZEVF
sBNUIiB6n4JiBKufaDjFwtKKKtK4nZgcnq73zbyV2y1bzlrj8yW1xwwseQTGlAcG2yF3ryqO/Nf/
A8PGqfzr+skoYWAVlwkOilj+V4Y/AjDQp4QfAwOkSB35AWQeE5ZcGPLKZIAJM7Lpco0hUuYGjYCb
SrZrn51oQ0TMMREmBy78CGQTCVNWGrkP0iaR+a4gPO77Huh4w2bhtbTXN3G9eTxchDu0WNKEuzSU
PZtgnrRwbUXzWEHjqQR87O3gK6DO3MlzuUnewL0R53tecJz1w3kDEh07p233PuZ/FMuPdG8khV07
KZEebn7IM6vTBQ9+qkzLbxpAxT+Lp5glCK9p0u1gIQNqeRyWKjjvdTJKhyW7AsHvVfLBH251Q0LP
GxlQ726Df8A7uDLfP9Tu25hUnTMjot5i9Kp3BrTRzmZcyn9tPmV4Snt3IGnkpdP6QVUZyrKtkN5b
hLB0QDavfhRk/g2/+brwSo0tzVV8d+vsGeDb5oYWh7HZATCBNo9S0hhYnTW9dRes7Mqm+7IZ7/ie
sBR0pPhqr+SLJ6T97e1eup4D2qIH+XkmFCuDCM7j+rlWgEwCNzlbbZeaxsQ7efx+OhwL6NwShaWG
zzW1z3G4+Dsjqm2zeSn/1CRAJHZuUcZUMwN1bPOpWl0q0/j53WF6j0qFj189siQqwWaSyvg1kMhz
tUFk1ouz4gJY95O90NCtN+32WpMlIFmQ3+V+b+e5yHi7lVn8YE5azNjBAdMceKMX1aGA5BIxaASg
lBdqsn4i8dPxAr6Hs8Sq72rVljQ1ZxOdUfXSEFHEnexLm17RsVlkP1gTy3pkpYHL5vY+lFB9GeSK
nJLjrJwcgLgBEIxoePuOkzANsBIXQ5KbNwuLbY1A6zu0UNQBRofzaLqHFftgVRxEKWC0+0Ny2Bhf
uUavk/wPx9E1s877CPYWDDLmUnVPzGHaQXL1x0Fhz79LwFkRq4q9HLSbOnyWx2+EprmlUP70zdxt
W7gd5W9HbJC53ZK6V3h43ZVaLDacFsfWMAXONURBzg8rEBPXo4uKTUwKrR15gVw/L1l1R7kia3IS
N6S83YuMgbCbm2dLlvHKG0Be1k86nGjuGnWVkjjSh5f/Bpwh/seoHCM0lKhGFRp4jNto5aAd7OFQ
Goew0RGG68Cmi8TB7ia38XdkQGPQ2bdYXMVyIU+0ESiGKwa3ILVx/VQd5cVi2sA/JKHa42hJ+ui+
HMhQdMO88fN9kMIAdIvZn6XqqU3tn3eKYMoBu7fyDMxL1AwtRdeDWEj6EuV65f0T7/eS2OHiiAqy
MGcaZ0KGG68G3yVMzDDaTOmNum9rOJKbT0vnm4SPZocelSNzkmJBD8TOzy1qFlilDLPw4gex/Loa
sEmsHIlkiFW+nl2P32wCoJs6VYhyE5lR4vOa1I1mqaZrarqKIujELJgYP0yRo64yfLu7wfPffiN8
EqMwVHTMF0yORyW9jQgQCNSulHvIzD9VfulRDR05nPUjBNUwTJXEAn1ef5PNXt9gnAhQHfYc58tD
N9PpdBG+7QhEb8WzrhjscEK30r+JpW/RjJRnzQl3tHlejyl+6qbXqBal1OBJMpeVBA7MTj5X9iRw
Jft2IViA6UOvdbhloGeR42q8kl9KBEaP8faS0kX7GIG9x7phR6UO2urh1QENRwLzq5r1bIWUHn6p
3n46ZWfyL109zQofXaRNg4GnGheycM5cVzegfiVPcXz814RsqRxau67BvVLVEPmPb/s9qQakbXVM
dOPLf5av+4Qe/ddTXBB08DjFfKqu5GQBzFgftJDu2zeKbuwrUXCBT4L387pgbVsHS21xDUWQO1IZ
l8L4vvgNvxJjVJKDjbjVTjG8qiKpppEqPTazYX1Dm3kB5wcUGeTdlcuiyPSwpwjR3p2Ql6tq6KM+
oSjJRIACtU8ywZgKh6oKqFjjY257TGHHB3BWJektuBCFgqybE7o86bHedLpO7NxjgyVy5BUJ2lvq
jA22Z9UOxwdNrmeXs5WARuPnK+VGaMw+ze5TLNIZ7++kuR6tcLZ+j0gte9Bg9WOxuJejdlnhCLWX
wdjB0FJT2OwD+fOO74/w202FMbBeHYmoHsoJ8VffEF62VG0GIt5msR8+5AVjUc3DntdBUHbEI4Al
1DmGxRtdRUxsQoBdhvDKbcyK9C2FvcaVO6igqzgka7XIJjcKIgIJO41l9ZgP9FsGMpBi5ZKg5D+o
1MiTEYLP0XHogTkDxR+1AjICX2rPUU4y5CdzUhpPPlJpVp1RpxvKJn35qfgUQLaaK5HNbUHC92LN
IEjkNI7UipZ7R9U2X+1S0t77eTQJgdhQ81ogOe9zX20AR8uhGLtgL8gpFFBqQJWLcOmipWthhfjQ
x9ByV3hqumfwkPSUL6VtTfXETM7J25FaNJLc9Yo7M0u4dUGFq8iDk7D6JahC+IEc8wsPSFLrcnkq
puWyFJ4nCMyC6ZCLqDcUyQN16VESqeUxvtO2vrQoTpnOQxus3Kifb4c/nHtvPs8SIPhWQLvg7Lu0
R14QJiMBez2pqIb7422obFZXWMv/3yZA+aYNULe72LeSlurwULyCll2qx+l89Q7HiMWE4/4ckxLd
WhP4galwNPmlFmWFZ6oxqzPzh2YxqC8WIRu1ZO5dj9YgGlacxyY3yY+BfMGJyYL0kG/7A7PJY7pY
CA/w5HQB46eQf4ckbfCk6+u8vq2e83AJk6yrxkikx+R4t5KEdAg+vsCO8jt0mZRNhSW2DEdq542G
LwKKwsxrqlb4r/t0TSA9Z0wrDdisTFVym4/OtPo4kzvV7RCI2H3lm6HhedNx22kicJ3QIWshuevO
pLVycT7Pr7sOUpSGIhk9LB6y7z/fKLfvCU1Ne1ynKEN+wCU3A1FR/MJKJtrf1ZDONnR2Hk7dujlC
KH9btJGN0x/6ZT5KjuFKr1uUZebHUjd38VJX+AzTXvLlXaInYkvVxSAdQiLlKX/Yj4zsmlDIWBly
Zok9rCeKEhXsyfsw2lGOHEDG68aSDCyUa7zgeRuAch8IYHWFM9gETEDRO3bX+siT2alE87+rVI7/
9ZtVKL2S+0POHximuKsJ626mUIJ6BrTxtV1NbhYTSw7TY+wn8bXldtRxQs26NyNXJYodwI9f/YdH
IkC8qMQW09qGvip/ZNdJTwv8hL5l4xOeDz66DIKFog9r8Ty4H/b0n15Z9k9GycqPMXJgSCM49mnO
SuESJgbfElL+rKQEEt+fP1iUzIDx8mXdW56aEpVTPdcNBSmwg0pTPwRHkPfJIMdUcnpDsFxy7PKu
5vMpf87ceQW5C+EcKCgRqd4Syh2tNYFxWFtt566IGm/wLBIVorPCdXo3rG5yM9q0VmRid7fC+MJI
QEBWtsCbYLpbx7g+Dv/6dUGwbjkfI6HgpqhJ5hPwU93UqJlG7ylUW/vC5x/pcWTrt9EVryathG1g
mExBf7s5QA7a5FfvRHR3dgJuYhIYoWEZYXrBoBEO9C9/I6gAEZRo266LBlBQHataYuWxi7NOgYjY
KQS7UztvWdajYtIT5MQjGiNsT8s3BA/etZ+U0wwklff++xZtITio13qaqfhLWpsUF/g01uE8Uwz4
+6Ntfi+Evgyx+WwZI0mwRIysSOfnCOY87P3ETI+ZfPJgGVoQNwD2GL1ODmi90+nkPLiF/hzHiB26
z071Mzwmgi+/QsJidurtCA+QKfK6NrPGGlk+2VdPPYlcPmoLuxbtTlAwHrKvBegzFrTPA9yQzYrw
taVa0Ru8qoWyWyx0mIr2X/YuLkJBphLXq5VknhaFelFPfv7FJ4bgFXiHHPDgp+6IgtVpC0YGfGzt
XrH29bQMrKiaV9r6pB3S+YSrcJ7ZlusOGUGFDj46YTy4LH2uKEsUJ1Yp7Pu0x4ynPovR1ixbK37A
RNAEmpE3/QgtPljxfb7FNOuwjSZC1LUhWcVnZbUeegXxFxRFfJwnKtSrjKpa0i3a5jue9g9i3xCu
jGFDVUiMqQbjNPoqz3pdaRx4rONzIwWJh2GJB/QbYn1BrEbvjR2fQK4PpE8iGs7Kw1bv4ITJ8E/h
3P0dGx+gH1w0SJwRtXyuMZaY5FTe5Gu554/MJbcJDWfTaAXSwGBI9nsrBkBz35F0hIHBMh3gdwr3
cLjR5JSPStnkHDwMyzIALjkGpoTAtV5YfiLE1YWCdrGtLvZL1k4qQwef0/GEY+FAG8124dmikyZE
X7LbGCf/AlgoURL2MUQPNfnEvZH3HgFYC7OLo9GkasT60i/mnmSYq54UoiQ4c7+/oyTjujOmMJj6
riOXiN2Wz56ERgyqNav2cI0YZFtfPmW6T+E6esTGj+fOfqiTX4eab75rSAVfC8Kqs7QkacAucFs4
XvzAH9pbTy6LZPNglVCtUlSBZSRJRsVkQgoajN1MApbeoYHsOSkF6cR3FVLtcGhL0FYkZb5u5sEJ
TfVkn9+SG7vU6qkAF43kpPC8C8t/WnpnjlmNuWmsGYoxZGo3nFtTpP0/4eUBDAIXdZCMQmb/Oyxb
drl2i7iul7IdkhBtyuGfvl3QdieC05nNhu4RWn7DHeEEAPTErAyVm033BxtBgLyTBt+mVs7N0DqN
wGgcx0T7o8hU7GHYIENdtORu9S12jd5yQQygVF3M/WwDb0AIP5QP4kht9Aso1tX5NLmlIlO1v3iK
dESZrBx5/YJ5+dHFW0y7Q7VR/JrEW0vjivwvQtHnE/LprhL1a1JqNOoS6fA8fQehkabLMqRMril5
zOAI9Rniaeg9J8rt0lUFVhWxrhkLUP1X14eqUH0PoTUXaqFpfCk+vhpasmkqKSTqqHrxrVpe4xkh
AFQhIqoNNyfevT089UI/CngOKc3YzboyZh/txTxePzw+bbnLqa4JaYpqMM1CFRvjSTcRE+mUernT
K8J1s/RsNlD/7YLNp3FfFs5ikLV+eK5qE59IYSGsoEGhqcn3imy0gOA+vAndJjNlxt25BSGRXYY/
Ctd3Mo60gBOO8bh7oYZcfLayHCm0kAJZ3/+IOfgdh6Z3VsZB9sn6kMAb4NvLzxS0+sxOHtPsoLDH
6jrgkqbhWQcFp0XnCxb+CJzxv8/kln/plDnLeOVLNrLrhYmgdCIXaEkEmEztNEvo+EwQWz5pDtsa
WLC0H7pqg89paU5/DmbsAU6lKxIg5JphhEzrSp5y8fh8E3JjeIyRb0hu5dW06EUVfEJQWfrXjL9q
Hc8AbuzniW8RSSBMA/Xns5EA3oHsijzS1CcoJTQa3NNTtvZWSqXl2bZy0USzw7r7LaftQ/iZnSjL
maxEOovW4jtCbPMG5+XANe9Sqyos4xxxma9R1sn+c2cudD9x0uANhXWMmHVr8SCmRxOe2xu/hFlO
UEDNqTJxTMSkN9ZD4PMceIn3TxY9DdrgEbhKBdX8T6A0yrrvfCcBltZLn47WKtG4amTKvZI6kOJf
tVJ/T8VEEa+fFELh1VBaN2Y0i+QIkPyMyKZ6Oa/zVscdKkZvkch4bIxAYTrfkIZOBcUGCP1vBYhz
InFunXrob/lbvWZWLJB3VofjUIJbsM8yQJUq1diLts8dtXni5Bsb6XFaeMc/pARNChwIYOHGtD/3
hxIIXidW2+1bb76Zywa30XHnzt+fyBLscRt+HKJkDy1qpaGAme42juNSC7eq51H2qO2kbOK0mLqK
TarRV3340asjOPI40tOYqP8qc6tBnZrv1KTDXeLk8TNaTVaPa5XkNzoPRmS5LoqTq27osogs4W7K
TsAAI8I6ROf00y4HDJuHs7L8692NtR2PZFBgAHwZkU4TO5cvAsGWIQQZdyUu2aHiDKHkWFeNOGac
T5K9NNkD4NQJ7QvYQnXLyUcWPiXE+Zc5aAPXtgNcRAgzWZqUkI9qD353Zk4DdG+qLGpKeqeCsazG
mK9uPl0XVCla8OURrG+gVuMasUx/Ugsbot1uaiskMNbTqFyKwmdohR+NhMsonpKrK+0VTh3ciLvJ
g3reClsn3nMjT1K0OQUnT7GyZ3WHm2E/9yqEcMGm6R9/OmwgThJaGxBuwBclnK50WMl6PAy1Qkt6
Fevdwqi+v0V04bJ47nIHztDP2wrkYRxAyXTYRUu+Gdn9renvC8mFtc0uJAp1CUCY1EHcxyblOr1r
/IHc3OdDMseSiTiCRP5ojIG10RXQvkcy5aswEzfbnpv5GAXLQVEL4kKac1fcDULX0ISylrYD+0mG
VrNJeVqgRxXMyVZKhMjnLWq+E/fBuO/8ORoToDuOeOP0W4LK3DdHjg8Cr7gLZ00/xxnwuk75GkEl
kI+12PkSjvUurd80FvJkHFert6RD/NCRjJZtJXKXRojUVzwk07/IexLn6BiADZKzQsc8JM4SonOO
69kzTSwGs23CkQZbrxI/HV/NDunaD4TvK7sSNt3hHUUtynVIVO2X3BPF7cttOIRrSmN3odQpv7gA
aRuKWFaPXF7XHw8q9hoG8bNZ215r/i6NHamiAMj2LFP84WW832zrMMXQDNo+SBV/fQTcaiquLVQz
4T8nRybSk7MADo6dsAvlel9Y4+53WWgGXucxZ5GyVUmvqcnExRhkmXd4l2acYQWQQjxufGX2OkE5
sKcZwIzP/uo8XWoRh/7bu7FhK4S7r43GNtbPwJI7HZnmRXe5b2Z7TJ2Xrt0zQYNR+2grhhywnu/V
uDFnkVeeuQMBO0rOCPnIoV7N685K019ynIYRiMp1zHr958QYaXgfMJK2cg/A9BGaCRLp92iRX4YM
uv6CJW5WLCYYKackoQaj91Uk4ogpCdK7kiuKKC6/aDH58DXII8sPWWRW9kiRXwwFuRoHUB8m12lY
jDdfVwxVusuj5QZO/gk2ruGXv57yPKLtrEAJVa5MFFp/R83/LYRJedWMkkIABzvlyu/ZpQyuI5zA
Bt6DQIRm5HEyEO1l4bfNGS097ZgSZ4yErfD/x/IEnl4CRvEC0GrYLSX/F1oB7G6S+VBFgiGmfHG7
/6XFbs3w80oWCqe3JIClerffDBFCO1aWn+bLeDn8Njao6ZyD8g5DqbXQ5wyv1JMXW/M4BRZo4mGb
sQsdMYPPrvEB1N5dZyHT2v+nrgMtNs6ngCovXDSjjAku4INTmdEQ2/7KLmGVqbqTL77g8HHhkb1Q
wu4qi63vz/vIZYmu9vqmRYOrWTgYBMXYe6BEuuYw6eLZv8esqfqM/A99HdTXYCWTZQo/9hDS5c3P
rfhaNX7Taz4/lN9WEwSaIH5tlsp1WcTjbjdHE/uy92+K5LDmU7ohvqJInyqDB5D88Q6YATRPflNk
X6xq1iQCatTOb4E+DxmWaCYJKn+fTvK26h411hfz87GMgYh52JKMIFNzn6x0M4AAAe0qLdxsWyef
MPumfcILJ+r+dOfZ9HREMbyg4Wi2Tthb8VEdDTkF6cZUKxgcV1/U1UXxFaJ0dqv7ZYzhjMsVmAGW
y1FpR3xZHx5Dc58McQj+c7kae6xQmuxEz6PQsGoSRTxdm8YIMki0DBhHp2n4BT76evr8VLpjIKIG
ydpb7bvZygpEAgGsmOlNduSyXMrB9sHZEBrOOKXd79pDsHrtOEi4uQvWyMlx45ynpJUKWEJjGvQD
ApZwC04QtpXo2wqWnTDg2G/kT0cBxh65chFO/uCWV59kzD1eTtHDC8jcxRL8Ep3aQITrHhCiLm/3
ipLG508SrjRL+ZaBTgBNVeI92PNIiUpDGZQJRDfEi4OeZrXIMrjRwg2n8wFd3mOSrtC7n6JPicqA
631Td5SmzSmF2pT4hHul6IW7bLCMqYQWFC1INKrWhk1QT2R+E3hNCopWaD+MkohN4iypTnZfxc3C
ItsTQcwE/1OhWAPuP04Ph6Ua9kCyQ4UHvizrrb+80kAHXpnnVmUxAEs4zS+uqy1UTiJi70sZZqfy
8rYIfJ1J+jvtUbAI2BNCzFTZMMrtJi2JFaiOUtblIEHO6hanU2Iop3OiJu1lEMbydUjeuJM74QSC
ap9x4ENVWhhbEKv8TO6uNWBzXOixpoGwkywPJ9OSDxwtP2dMRv1HEAjnTUwSyjO+Yu+Dlna1aFXW
mESVJ2QNMSF7818tBnlLmJCj8oTA6cDXswtsb/9ZRKyA6WDoaY+JXTIFQPOG+rP/7y5IZitZ1rK6
AZCvl6Y18P72MefnpGnw5LsNRlf2YEyygRzOOG86L8EwGa+lNyo4LlR0DYx28y/mlc5nEKxHekJF
tz8noAz/IF9bJJ7J37Tas8LwHthJYGypPDmxvrPaSHvjs1WhHk8uwfx5EpCsNFoqnUXsmKteHod9
inVa+6j5XVePnNzF7Z4R9LrQuN6XKDzp/tSk/YL/x1YGyUD4d5dSNRK0/VhniEfb7GGSNhPoSK7Y
48zJmmaR4IwIFrhAi7yBuNmrgt49i7NBzM1su8yaF+szcjcsd0bpjC43S0Y1oYrC4KDOcjf1x1AF
Dhu6+r7TWlw9YsrcZKvE6roXvi7UqHnlJUjQguEgzwzOOOhvmkQ6185b7T9+HKDKlliAJPomZOy/
jXvuLJh1gf21EoZsZaH6KCpAXJw0fc7rS8uu/5iA75LJBftjT2qlSw/AxpFePK3wyuD7pNcFu29L
iESuNpXgjl0MYg6m0PbO4DE1s+HeN7P/tXGNGjOApKEtgI03AVFQZ6fkih7HSGAyKq7nDOYw6jtz
urbMbC41gR+EEdbpc/TtBCMRNo1hOBHE+RiXUh0DBfI049EnI8+/Exd7zdCGwx5wZoEps53LItsT
Ok05pt9I6x5lkpH1AGd6weUFVSONZ+1bIxi+ii/3Cnwk3gk0Bcx+w+jWCEIs5WfZTCMUbQhupKUi
IZUsiMudDCleF2FJzNZ08q7oNO3rgQhhS6QnCABgFS1je2fbkIwgo39PyqTq20pNU9ObNmwnsR0X
K5nCwfNWyRurXdfxkZk58qDfD9ud8H0T8igxM7g1pX5oqBAuDowCzKhE0Tk4SRpru0L0e4o+sEA2
aXOP0oxYqZ6Sw7Gws52fTGr6gEVeeOfDhvsVX+hxI3AYnmc6UtFETldG7C6kaOzCNo/9fPxreh5i
HzbMJ9TlSXmz7qXPeidm5IExHoRIdYHPjWC09eLzJkPb50VC1h2MCbLIQuHDa+82geMbPdvwYA26
6wRyPalkYmiyKRo9e39KcFN38FujR+LUc5Qwoi9Go05fEhvda0Oc/vaEqSGaloAkTiHSwlEVpZo4
kN1Pl+uDHoZYOxL7/NGdYMy76gOpbPo9lOP5JlUAt6HomnW4YoF7g76cN+z4D/EEZm6CCBTwGPYP
dJJo80wbfy/EyLAru6Y+4cPHO5z4e8jkXkhxqpXAlEjoUE/dN8P2yK5SJFK6T0bYwTuN9QvmObTY
46WArV/0RKjvdDaH9TVza9hcYOZHE9YEgv5qubRiEK+kYu/oUfCWZDHIDjSvGZBrLqCE3gyobS/c
jpmEu32wrINJSWY7is5vcUmibH98Tf+2Lq+eIrz82CH4wG0t8fBj/x3jsDProrpV9KS+FXwSe7P3
GuaOG2NIv3AsWny8CS0zcd0YFCAUdhEfucPJ88+zfmmp2pGWXn8iA+a1ayKf3vQl8N6a8hfNjBJ7
/7vpOhJ8/fFqdwlFkeSK48tpTRyWBcUMLxw3PTd//RDj+CD/XhIHlDR9iEe+aUiAKwZqcMtlsOJJ
Le296D9l3nuqzrCqgnRcYEQgdOKBvWVX4JsiVoEPEJ9333zjRufdx9i6sR8aCUGg8s4pJH9DROPr
WO814A7Y/usTeS7e718g7KTtOiz8dSM2zq1m3CdHJ/nQbk7RGz7TMgQlskt84KtXBsij1HkPXZRr
QgjJmwY+CSe8KD4051p1lt0HHUmP87T4RGjl3qe2nlDRUGk/7S1YQD8JJ7tAavo1D992g7Evr1Co
DsMhZyyjEZpt6Db+WSmLWKF7ekF/LBLtMnYf9wny3cQtflJOcQAf4Ic7nGfsAUvbGNu8vz+uJySI
8hCA44UFe8UhCF1b90LUiRe71LoTV49YXs2PEicmIATfnYON2TMSX2rlO54Kc3UrmwmJ6rO64ux+
fR1FKV8ofGxdj9mOMOIm+UNWWOA6dtqDsjY0CyYtoo4364Vxtjf0cxRiFFka8nlXHNAs5wSnaFPP
0R/ppeDDh2gXR4WMKXLDnGnUHmh67RSBHZ8ZqapsniB9NJzFO5i1vyxS8omixqy/g8KxfNjaiH8N
pE4xOoyIFOjA3Rnx05BefufuhpNg7BqjlZt/1YwaUyH7eyB4lVq8N95hMt0m94uU69ZIY4DgLLDw
dGYRVVCfCYieZSsrEcnn48i5eukePqIrW7wZx4TJzcxHh+Eo319U40qoYrkkiGaXuIJA6cxUMDjm
zEC4ZnwtdIX8qsFb0X8xDhnGc/uENvsATqIdsxDN04lqSegNnikGrwche8lYaoQl7ix2oTo2Wb0i
j8mSU7Uh+WDuNSWp8e99tc5pZK8SxO7k4ry42HRKBUc0GaJHa8XKx14fIdvWegvd0rnrOJDIJGH8
nzeqLewvxNWxrJYRMEAphdix07QuSlApHOPYDD1NviZSPVuProYYiWccyQFi0NHCTvuiTuIsu+i9
kdsqZ2aNeoYQdLZCIPj9U4fBagHA1obwNALYlSglGgaGTfoZSkxbt+c+MaoHxQCAv7Hqiznr7Lhz
UyDxaMANkiG/ZhwyflN9T438RGTqGQO8wVeqh1hKjR9baDEb2Exa+6wbaZr2Sql9SIg3qu+Ofa65
kRcjJ7b7XCgU65TyA+elYqik/FExiliZq85fDBAo461vxVZ03bYp+TbzsnxYEeJ5PHiUhncA013H
Wivd8tvM7jEwYIyF7zEZgRWPbWE14CX0TT0oi69A6LizpftG5hzJBrphBMsmKRxh1fny8ccWlT1Y
+Y/NeghXtvINXqNBa1RvjUlgjAEkewJ7ytJx3m0pbx4g+9l0SU6d62yrvR2v4BDnmrOkEteifxx0
CR2ScAQ2bcJ20i9S0FSCbATjjype+w0yaCuhCkH4ypviKXNW14XXGlBL9oaDzpn/hddXw0zQZeOb
r4JDWEVvZpUXd0tscjexrem1Z8a0cxgi9pZ9359UmqwtTPDflDiYnQ8AXIib8gcaF8nK6BKrBi1/
/ZzrGbCTfncRJ2YeZrz9vDmXUF0Gp18C0zea4+vfLbdAVeSeoqNzLgFqDpg0FgVDK502KqgCKs6a
NHUx7DsSaJFZqjkjbxdc6yOSrsIpDw3UQJksBEMHMNn/O5vyhdeaxn3OuHX9EVZgXUEsho0IpCv3
Te1+Jw34x6Nam0aCs5pd3uJe4Z/VCgd4TL77MiQy/+fqrh7UdVRDszr4QCcaRetmY8KDSTJU7elE
Y421mGCdQpy9uVdlKmJ9FOBDp4JAwmNAu9pOPM/ybVjGHNjKmD3DTLVC274t/BByvvPTRzFOnWDO
ejYMVzU3LRRGJ/eNNrzxycrhFWsc/MY/EC8TOyYtliVM42b0r1MQpXUYUu1Nfmh8A1/kZgI9T+QI
k8Olqcx9fevQRPRIT7PAeaA6yqv8eb7S3dWCwUAtr11+An8HJoSGGGQmYQL7I3grHbPzdp4vbF7B
56ljCaTrukCYHdy/HBSVg6YscKVZ4c4hB7ahe0HU/7SEqg2K1B8SblkIpvIdFYr2vujCtsI06q7H
IOxv3DCJ+VelUkp0mcdOVD1ob3XXf4OMGBGtLLK5zbYHIohkJT5eKkeZXT5FF5kEwxavWalPqzhe
CC+E4WftBT0Wuggohd7pNp+q8SS/Is8OBz7Ng1YQ8c/I/Bg9UPinKkqfwkf7ZxOabUW3sXl7vHoV
MJq8mLZpi9q7l1BU7SM9qCYvIxqskr6IbcX1HKkplFdm9c+BPIO8rz4O47KYXmMgin7fkM9BYPf2
yajDFJcXCZ90nvI5PxXIYAfjUnCzeZ5f3HYTRkN5QnS9cOsnskpfGn3zuGhyQDJWMWx4FEKd7dbK
7XYEjq9gV9PK2xae1eN4L0IbhGsTa+H1XBhB3r2simkVIOKjP44co0SVM6wR6k+crGZUvInIo9tw
d3rHQPlu8fpyv5DC5rBapETt9sJC2Vjb702SVsUedEGVT8Vg+rqzarWma5QURk+2++qHeBjtWPj5
5KpHQiLu7EY7dD0bDFBML/eF8uk3a2eNwxjljFKAlA+NeKeFsSykp7T83g1YCvSw5+US6QXUu48M
o6RB3z4WGZDmZYBfIf/lMtDXMaFIerreOEJmNCEjAm88TfQyieMQvd5KiVcbxpB1pOLJ+Opq5nx1
Hlny0LecBJ8T8BHZBj6XZJ/Ezv8KNUsFlol2gM9yLRwCA7/RFs9JjnJs+Bux9q2zWdTIeWT7op/+
p2dvpC+PBzY0cLaA727K2SMo1rco8sONKxPy0eyBcnnxLCPKBpCFpd6H4QDg5CmsUVvz8k5oy8LL
XuWX6n2kpM6cT2yoJKKXYG5uIYLZrDYGwitQD9Hfrd8xEKSSRJ68j4psGHy+hzEqd1HUZSAl5GJQ
DPDvACqvElpYx1ZshyWGYF5ZJBTSDWpNC8c4NlsnrLtX5NS0Fv30VWD8yTtItTh/E8piszcrmyWQ
5+065LK6/0PRuqzvjb3Etn07Q7ChzbNPXVJ82cAxPSb1x9tu8iPU6kgNA4pdv+XDlBhY75XnkEqx
H0hcEl449DC9goSaz7/0gHF3a0Gt9xH8hH48eZPxfgk25X+PbnLPRnT4Tdu+Nu397kSoN2wvWG7s
wXNojnZlHIwg7Gtnd08qWw+40orLj1lp66H4j0hRr7HSkRfL+ASDx3yppm+sRTn6ksX1qUTDIs2n
6DHz8/3aAVyzUaNrS5t8arNHgMSAJ7RyRbF9yL5ufgEm04vHxM1+9Q8ueyw7jEfGK9oW/2CdKHzi
lJ59OK5PMNi8Sr45xRY8oF0HHJ1lqU9+WQHB2LyVeNyqwDoB/sttiUoMSP33MLEGWKqB02TSha7T
D3vDrKiJTax87rrW8+SuOI5AlRpdlSoCVoLLf1kqNa4214IIK1vf7Lv2k/6wcIe0vn1ZribTI0XS
sCg0ZiuHBId0tclREU/6tfw4vMlKQoA9+jejSt1o0BghuN77Yz2M0bDS6Y6CmvzxQMSFJtcTJ8TI
HjHOrLFlpMEnRnX+nbvKRik/vQ7e606nW4hLLN92qJ1ie5tSJNoEWv1m7kaubgG+XicFS/sc7yZY
U8ZbzGAfL45B0PZh6EsByxSwEWY6WIcJM1fnE/bTT+XgTbCEQCwUnmUJqy6jsZNVkCGUTMkoj6JU
qouaMDuTt8oJesyYTTwNytjbwzbYV8HlCPJhVWEwEWXXaBpyA0Xr4D4MCeEhQRVhg22vKft6RjnD
sE+R2DusQAfpZ15kT4y5klb4B91xlaZvvlBIN1keklcTMbk6YDg9w5KkMb637Sume3M8p/uvupcw
uk4mBnVMwgIMI6DdJ0Kc5JR8U3za7XEDIsMui3uQIWTuDSGDxahPFaEhr+0FzCrtPYXKvTxSLY9G
FTIGVXSg4Vs5FPVqQHer2X6HoyA3Im5NoMRDnd/TzABALnBPGm0MKufBTzL64++69VVpwisf7DwJ
xxVDD1QNuhpbjjxWlzd0ZvfXVqGCEpQhA/3Kom95ytNo2xeeNUm0BF4fOPbt9slz1sD15Dr56jPl
wHhq9yxMiSLyUlzbGvwqfZ5NqyN238JYV8HY5R40jGGpCM4fvcYfS19Ftj8o5mZp7iU2xDC7o/mr
37jOm1x8W+DnuB+qMsCRHf270xSTdNMDJJEZTTt3g4d96nfHSwyZaNCdNf8x4L2ULnR21K26NWDy
+nz4DB0zsxnD/L4rvlsUH3T13llNONqjcx2tk5YSp6D/rH5QhWnFJgDhBkkwEbiAmJKIs8scbIsk
ru5ucG7ow1n52FLN3zuZ06yayHTchMxQoyZ9pGIn7UzRSZ/0burJ62Tevv4aJ41wxwndG3/qLHEJ
VnDLER/676/DWFsx91m+pPwF6QRRm8lYD2yAP3EmnaZvLcnAMQd92m0G2VwHALyJllVIkhQc3tMO
R82aV5h+M3QfPrk9UFPWadWjDJSQBn9llNIeYbdWzmMYMuUoucqJabLwR1IuepqCePvbMie8KT+e
4vKaU/cgkWOWumsgm5rw+CDQPWK+EGHsIC8jOfzvjeAU/dZQ9mJvCaPwkErUM8ech1ECo4k/oGEd
+kTTsbGaH9w7D/eNVYJpE+KnwdyL2CC+j3Z8xU5om0YYI1iwlU8ugG6nVwB70+Y6iGi6tENrQxIs
JTmOsZdfL8lzxh+X+BvY/BhiPTofeqjVAa8kBKaP4lp110cY3t+6EhjlB1go9IOFd/AieVZDlrsJ
7C5qPabeBSWXzLA8+CwaXX5XIaTslpDtuXmusin89RZFfKlAM+ixoQyeAxGp00QoIYfy46ikWueS
4gP16cr9PXR2BnE9H7IemnWl7Ndo3AxefihVvHr0f2H9q0GDT1i5bMxhE1I3yDL5o3AmTlvOQ5+u
z1A0kMsXazDLro0ha3od3St3LT4WiBjLyWdlNIL9YUsEMw7Z8QJUtqCxneU523Mo+unclLPLt0VT
5kb9dAcDoCxKXK8sanu/KATeDzflDIyO/2BBXGv3ccS+f/stKkRhsRb2fVXIkSQQOg9T8i8bBJji
HnDNzgdqJLfWOFKdh0DwJrkwzxPZMq/rjH4hJlzldRmQ9HkwwbAHYMM3n64zLdzSguRCv5woGIJc
F9+f1UArwkEmVxuMD2RhALwpFGZRYmigbo8X05UsfZS5Dhix5bEj6EWw4RkqD2DTY7imt2nFHThR
/u3IZO2FhhBeKRRlYlBXfmWCI6xbj/aGttyqSe3Z0XaQKTQRkTps36mlijKvM4fB/U4vZkUwvhAV
Qgc3I8acoRfnQZ7bdSSFEzP1lVSH0DYwM4kLj4rXuR7791C7ZQuosYXgRkHBrlwyLimV8zFbSel/
ZoMgJo95rdy36tyUx+AVMLRUe+Djt8CJshtsv1D9nHTzaq5DOpLKLQ5A909N8Gy0so76Wl1/BAUD
b1AK/yUntOHn08XNRMsQiDhuM7Fu1jw9X04CbAPJq/tYy6+aQ854r6N6CVNIAggEJRvs8cdsRSyR
PaIpmSO0DMu37/DP9QmeHKwOCE3tJ+cSioodAstDKSNaO51QiqPQb4n/ljLMmli2dCKndadzhMeQ
h0Q/4HK0cTBANqhyPWdLplfZpPnFP3QidT4WBe8iGUd7Xi0dDdmbtd31vUF08+Ze5Pr81RPMhKGA
stNaiby9n+PZsGMnipxpyObqNue9tSYQfzHgZQEXWwpyWsQ6PIuWOV5WnVYnPfRWOepTYZNrnknX
pRS28RZ3WeSEnl3zIepth9GwZoX950M7aU6ss7B++zCxW8BixGUH47KQ/BmhFIhuzmsEkiI0fu5q
UeWVt7DGNO87hnsJbuhqfvrbKwcHJfAvdzP4ZYjYzW3jUaZ3qf46q1ghOgYOO2M39NpNtFXXvqJy
BmcQ1rBJ5h1Ly5NXrgLqNl+XNCevSarFIjf1J0ThoxWNRS5E+LR5KIF2uChjKnHmPBD0NJzjI/ql
PS9sLTns9Lo2h8ATbNJSc0dZB7Ca2SOI72c8mMGLXOYF/vtTcXaOdb8x81lGKaaFe2p6eHxLnJSm
r9rTfo0caKyRbB2f1JUU+qZ7aSFLB46w/fyfBYgULJM+gsy7cbpt3ChIgNQuArwE1Yc0kacYpaDe
U103tL5BDtJ83XDRhD7qlu5+vaM5GpzGlB4Vj7xAfDxSJKqSz2eqiGo7NMVgYUyC5kBMtecgQkV3
zD7HOhH9pLmIRzWFg27sHxGfIh7fbaGQnASUCDLBOm2Ws0TEBsa+2pk9bIPmZjC37WFsUBbvr+wg
jdkHNkCmBiCNSt2PZSEZdbOxCIjt9NGalddIFEOCZ4edQK8fW60BJV0RnCDWLWs8cS4R0WcAOzjA
wyoggQcAHGKCBtKJgjXC6EgzEIHcnUDhLN6hBktjMj0+4LtP5AdnMxIQ6/2w/JT4sgtECQhbC4O1
ZazwN8K57ACE5Rrn0xI6d1lYT7EVo5OnFBJQVZ1GWg+O+TqeDyjiscUrb/6OK11v2zQ7kEzprfaa
/ltyDhUZTKsZEfB2VoUEDiB7MvQy70Dq1rXOEUgjsfZsEbJrN2oadOp3++FnDR2XJ1lam67/Wn3X
60u+u2FyONAdnOa79Fo5bdkxwzS68pwZ5MzHEDOuSEmffn7PsL++pFJaut4EeurhU+HSHHciYiqw
ejxMJKVXD1Uzymf3ltZ/EAtkY1/miUCaghFcjnWDNV09XLeIEQhYF7Y5k7w2Nwu9MKFpOAR0VAo8
9xM3tAxCh2TlWJk6YXI+jUpJJkLi6H4E9/K6mtEMifqOuW8EUnf/hPP0vQM/OLAOgQJ1ecLYq/h0
LidfxN8cst6SWoATeKsFXnaeHRlTroul6grf6PofqHdF6Al6AX/0INxVcCRNg2dTY1qB7jTQi+2e
18IEOV529uKFesDnLVxrEoTxLk7cWlpSXKLa2JY8ke30BtASxhkmxnuy/SM5bWjKYPtMl4cvTRT/
CDAbYjVczBQmoFEcvjxuoX944TUDG+82choWF02DxDi9PVQfd3WyBLD67zOjtTzzBgkper3/hH88
ZvJisxrPMIAj1PVtXqhYtreVSSfbiI4Ht5xqDmC+iBwgm9yG2LiGDgBXgsvSyGmdFUxIQI2PV84P
pPzy/FyM+t8xMnPCI/GR3MtyNgOMIML04y7RBjVNsUamFAung0cYENGRfRV9W9vbr9omtYC9KHV4
jDewB2lOL/t7488oWSrWiHoRjFh/J7/U2I2QNhr4zOaTayv+KHLv9izTYt46a+4hS+VtzCM6yahZ
5N5IvN283WTcJeqcnPaEVhfzovMeqKPp23XldBj3lI+mFitHJGEuen6TAUqLEqHlDMia9C7rZRCG
MEUtJy0oaHzHUU+Z0ymYlVypuUGiDgpEwIvL3GXj284UOYCZ4B0MBq1PPm1Bxfa6twDOK3huZRAM
HUVuXSXF0O9h2AjF8JEamkwle93lXLubD7IA8kls/eXGDcDvbqoKfn0IH8J2DQLsrdAQJ9C/f9zB
ToBQycaMsvxlQaBK4y0BxFIDdHlMVi+NI9mmK3PyAMKuWyi7cuFOEG+ffBfNtE6DpieCQCBrEwXt
rIZLjFbulCa5wOXuK4jM3d1udJMrKfsjU5loZqWvZV6C+5geShA+Qqc1iUvDcqdsLroH+kmNL1IW
uoh8U3h2YnZ8275riO0sED/UKOzxxc5GvdIpzQfxe1oryJUXmaLIaDtgqtPJ5pO/asjcAnIWyStu
nkc38pdv/qtwjUxOP2mOdT3wNwjekeiLc1kCp1ox90mq5Jw8Sw7xMSSFSfOVL3+4jOXIVPDkEcR4
glTp/x6jweXb9+nIECkmSgHkuueU/wHVDwsayHIVOETemG2egTNZk1iD9ILmTUicOBZJuo+2z5Zk
D4Sa3BCfWZCpRH5PPa1twtxVLNZll8ayjKeqPDpjJ5P2iAy5yK7HjxQYTIVNPYnL2m6gDpUhqhmi
v7XDEXoQfru7RuCsIUcVazRpreCnZ+VeiFsMeg3aXI+if+cpEX/sacmEq/gpHKVszpW/j6hJ411a
xD10lB+VeHZID2gX5xJi0Nt4DaCJToD0ASTKF7MarBSyOZzmIDKYXmyyzrT5nrQAmSJcvzqMCW0t
FEK4uASZeI/c2Dgypzwzxf64ta8ZUsuSCoxAn+Sga9HMDHBWSt5g3u3mSdF3JWlak9Oa6gIXch22
LlW+E8bayDOQUF2/JQINdf8jW67ilDNZO++Pujzwiv24lwljc5/8+rT3ZBARrJvwh7ACtlI4RO43
uG0eAX0ULSGdB9FtiB2gebZhmaGcA5Aa3wihZC3/LTswycDOl5SNrV6AdcMDRM6XZzY23UZq3Ysj
IP9aMjIITbzosLCLgpcp3Gc/ESccp67txbObcwEUu2azscPDXr30b6T+KuofcRZJiPiMq5jEwGqx
JhiZGXrjpwaz+QAJZdf63OW046k6vG2Zq4xEyB8y3jPxOOo83yPB6aRyM9lp9Znt1wX3TohvKD4K
JQmX1lGginXfdTxpDxg2epkzCC+lDGZRLNG2foGAhad6+LL4w4NFnoGFpKbz+NWQ+OvIMELeIe1y
RPBjBP61bKyfRh7WnmOrtVOIA6UBzwkhwFcK6D3Xe9hjZIAr4DmJ3Ia6VnxR2RoJ+odOuErguEkO
2x5xMGa2FJkUiG7C32zzhfTyvejl/1uGOcA0cvSzgXlYAjZehxlhg2IIBJb2+UDZijoNJTX6IpVl
vSmfW2BsIj5ullgJ54mNP1Ygp+R+1uWK9hfgORw1Vxg2JixI7xvEVlwYWgHUeAItjqithlZK1hhn
BlZkua0Z6JDTbjZmfTpHthEvy7/JMJNT1WFrvzT6hkaiaO4ennKlGL2DagNUoRV0mo5H9rG1t9ih
4RcB0mLNnIVy8yMR0N4ZUft04W6hxtQ7zQjNZHOBm4IGzJ8Nxd550fgHFgiXLQAnfRJdL8IuVs9i
2dl+BKDO/kD0e0pbbrAZCcQIjknmcQ9Hele8JpxwoAnpE14TrkaPqx8FgUIazCed/a9/VO9KW8Jz
CVowmyk5+06zXf5csDCb6CfX95s9XnopqBdDxyRjg/64J1LP4Jt7siKAW3bvwobGg5+82IBhmdcZ
QkB/X/jR9cbhqd3Fyl/8XA+ksLkhCL2pcMmiF679n7irn0yDtdpmLhyQLsj//j4Rxujw798ein84
ZAcHVxf7YYMJcSyyW3P15IAKB1Gku1mPFumXm5HggEPyDUC3rVlT8bfGAkIa0hBHz9yt0mJhoh90
96tl3sABgCEhwEEJS8nLqOIqbC0G0c0vzuKweRAygVkaL9tJBFtdckXgJupYvXmyo1r13slIT5q8
NGa0nx+sJ3L4+Y1JfGxN7KOpIGvvu65hBVbtDTHB5JUAa6DouaNbDbQiCFWwuKz2i2SKyVAoieaK
Ja0YU2A1qjiQp6xQUVwEi+ZagoMraHNKf3i1tQEM2RpbqtMT9pgi36F0pkLdWo3OfygtBXdrfRE8
KDEhUGx90AA43KbF98f5L7Fa7WvZPQEmRf7K7GL2If2aSQgkH85q8xi3APVHRVdEu+2s59jKzXft
uqYClEQoVA3SzvtlNCfY4wkmJhuoE800TMQfD0k7dMm5BblSxbPbgMBKf09dHIBL/zj+mxaghpu3
MjgvnmL5Li6/lQwfFS5neK3/GiELxN260Y1RdwHJ+CCVrO08LCcXcnJ6vBPirzR/zlmy6IkUtJyl
Zsd6rgtEckkZT6/mjADBY6GfgOJLO6M07cNBcl0egIn2VJJx5OLvMCtpSF5ipQhR9JEKdv609mTh
mU2jpIg1mhvJ/HBF4IgcphtUIHLj96GZTlt1WErR5YHlqOKfsSpZv6toekiHjq9giA1c4xXQmfUy
1Dlb5G6RkKu5nLzxJqMP+2gMV4AZ1/tz1vJh+fqajMHGYp0R9ihIRYm/G7jz/41ABBmUp6p/HgqP
JXwBizhYOAsL4VMPDCrT6TZ/tAvgEIecAlWWyZc57GhBbMtXbwcjxOoY4ab0SBIb4oJ777J3WDlt
VhdH/HVDT6O7lCtnugrTQeXPOU+4aWtGvV1Wk8DeSJ4GOyznGgBB6E/0M89iFjuhj7V+1R/EZ2Tg
QCdT2HH9WglvzqcA04juuFHpnzg801++k4RW+Vlks5vKxtpEPYZovaqhK+1mktJkj438jWI0VHbX
R1++kZN3SPJmzcG5h6D914XV0osNd1GrKpOw2CXQ3fBlD70Lg7bOmcj3N6ZskNoc7y5Y35GfYx8a
l8g7fRLbWqj4aHdMA6hwBzKyNRFmNObGo+kE3IkTCADQFk9j+Go8CLi1zbhNYNSngQplgLFE1LFi
OaimFSLErUCkG9fRho0cH8V09EIcYLdmmG9gyiJVmSp/ZhIwQAWAWWoqDfmmZUzLRunNfZyUXbBS
NQTxIgbjPelaGs3tbYr5TNex4QV2bF/zNsKpYOMJg5rdWAm/EPyWrv+w4gcZljcoR56dtp5Ai98O
ALmmLnUr32fWrvzFSyIoTGCOhrgeZKVsmltD4A5BxKkWWWqsGcmhQYvSSgT5k1h0aL97etFUmpGl
eNZniE61dloOXcooKb8ELgf5txpyjINMQtpsdTptZ+2vdp4y45PYTr/rRQ3QJidosH2V4B2t3qHP
3KGhZZMEKjzSBfYZuOeuc+BT3vmt1Fqrxy7C7sFm0gdDhkeSFem9I04B3sHN3yoaSFHnAjLEHlxX
fiSZ/Wu19v7aVfnnra0zBoZ+3aIqOvwrbvXo/GJB7W1vPsoTPgJxAAhndSqhbJuj9d5i5PKeESdx
UEJM0VvF2ogwp+jzqUHHiyv0NuEg5GNgrdcciijR7FvLVe9n+1Q63U3ogoQqIhD+PJCxrDNzz/R1
asLzZce7InfmmGpY6EGEWPWyxui/qAj73aJ1D8rfPcrphmSwoZPa+MprSvZtHoL5L/dKbn6UQtZo
WW+yr+PPtblqjJhbYD3R4iLkE7RhUVR9+X031s6eYFA9Oa6nzau7Q2C3G32/fx0ysMZUhiV2Kb7U
m9G4tjqdMoq1mmX4v1lOMrEdSpBtKhIETqBE1yonRKyz38YlxX7fiyXAs/LUzzliQSb1ZUarw0mU
Z5w/srZ+DLLKEPQ4dK4kMFNa0g2uzXf7DmFNmlzOGO9iEafsRDWvYnAwSuF9J5RBQ4Y27BBOjo6Z
vXq5Bbgx5LvzZeP1G2TjCSxE78NRC1CXWWVPsqEna52YELT6hwNepHF2CIySmbI/GX/YTtiPqZko
dTpC1Ro831qcXYtzJME/jwAPqd+4naGU1/ifFAXJ4qnIii6f83yIGrvdRCh+i4eRndUOXbUyYRBD
LnZg5ggsDjU76Rd3jWQWWqMJzJ//9Wz+l8+6Yru0LOMWkXMcroWa6JQ445fNvUv8ePD1D01JYQph
Tna/0nWEO1azjtVukwy57UCOqP0HO+PeGt3nENvFIdqHtNwY0ulRYMKnwGqiCoOotKkgWwl8PFct
RJoSb2IrvN3HqyUTn7kpjUh4vPBf9EbwIhgXWtebUwg1xKmXmpAge6vEFMSNinPw3RiabWs0xIFZ
nL/cH8CvSltQG1fG7/9oPSsmHRg4J/KPhL2gssUaa7QY0MCT2zmqMUMmcVvAF0jg6jt/cG0QjKqE
yBQw3bC217ILUPtzG5xkU36ltNPmGpnM/7UJaCg3BGW253YWZHkLeZQNd1HXANtt912ZbT0MV2sP
+pD7E9Ly/lzL53Nd50SR9c3u+LN/69y0oKXM14wMD07pZLAKgdUPzKZzmVojAAM1r4z35K9hj8F0
u0VYWMFjSfd/yMS7r5Qszu1d6k+oKKAwxh8tGF1Lc6NNuj1ZSOqcRHzCJJ7CqCwqqbQ4bTLve+JZ
uMmgNFnyo8HUiy18rLiTLTmA+dvqABV1GH9FTi/0HSQJuy/NPFn2gPfLLrEKZxZD8m6nGnvhG738
sR+dXz1bPy7NYeoJGq97Lrstz4flcNOdF2wJydxpPck8TL2St5MFBv4XIdT12E1LY+ABrzhOcbw/
4CWTPucCeHwg7kpiJIH1hRnnd+wkGFr0zVkULZZfqbG/jXg0tYS7agH9MlhyLQ3PNOexvnxSO9fs
tUO3zl3rVuJO7J3xnBF6Pdo5SJt8O0qL3TahJoJtWxy+lMXKnaD6LcMOkaSHDN5LiL3OVjZoGgqc
5Up9DKJ7CH5rm9wC7VoPHnbmzFDal0bs2SmDK6w8Cy+sGrySSk7PcLdb1bnmX94i/Z+us65yYIWr
LyAd6QBN+28ewDThFwd3h67xLSA3clTXR6BHxXRToFKihUdrYfU6burzmyZe0xf2JdafzXzyVp/P
XMZwuBuu70vxiHAZELkRQXLS3dkNcjQEy+XfAXCGhr1g22jYALtUsZqdTAPVBmx1fty3T8rZFtbO
IlVipM3iBL18PgjXZGm9UZHXfT8pkyN4N21WvtYtxG9s4+ASO+AHTcVPViRTvtavR3R9hseIwVQ7
aP4+GjThRP4vuYP8waGoTHwn+jLaxQf5R+03fZEyHZ7PKubuuO0nD3TBBSdAyA6m+DUP7cwVmYbK
1nNE9rSOXNccfbb1d27Da0IhzD0c57GgWTslUt3uKcrsgOje5mIoE8AStsPNE37uJ2iWH9nyHM3/
VJju81u8Ybj1St/LMMv1DcuOZeDpu/kyHog+Rs6jeyqUlOXMYjub6mQz9T6HBlzCzSDUyZ/8VXTE
lHHDzuaKZzrj/dw5XfYtXaq51n3jUYBQ+NAqqAJJiDcP0X86qROgXeBXUKbqM1WxDvZ5/2Jdt8B2
YmmzIN9b2iqA/wZe+fyVdZxbXjZdNWgFxE0ELKyleBMb6VUTnenwO3/6kDfSB14+ofsOo6fQJGh1
dYiZcCO6gcolbgYjLbQvAyze1/VSM0tsdcy8R1DSkI1yqQ/sjRIS0PI0qcLfIQ8EF6+5W7Dgb7Gj
j10mHH3QWQNTMQju3Wlp4atjLfJR7SPZEbS2kT2ooI+32N9kgC2NVzhEeIfqV3JZ6eH986EJaNTV
K1LMyV2c4FNdFhdIoRobUc8QGR3H/417tld/CP1W5df7SlDe3fw/bxieYU3iV7StRwcSrdg/lxOD
4JlWXMuPfa2hNMnxaayyYfT3wCHZ7ueUwEouD7QpUyTW8TOdcY6mNv9DhkpJZ6GJUjkpaIok6Oui
Ol1vZ8dMCogeYDzvJFtnB/8aD9dUa87eJUVn49j2umAnbJxQRYNXaqN7f9QoGjcTfVeiBGq85Kxi
rIEUvB6nToPZQi3TBIkwo/MLvPIDYgreVyAgT5YcHvnctgA/tw9pi15A5uAxHxn9YyF5gmuB5Bvu
0hBnKfp6NBgFz/FSWTekPjdkhMCt/VXsnFVGS6CkjsuqJCpLU82yGIYIkb8zhBr8nWDmlG70V9SQ
qAY1iSLTtLp0srapMetfERo5IP5dQZSmG6/jyYdufU5xaO+FC3Ycu8rdMBmUYuC1PNjS+pqRBfRK
MUz7LhlAYHTmBOmkDhnox0vZc09l5OzmmQ2hN+hQdVDlpZ5V1pmlQZKUfCPN/ymqvcAv1hUjoVKe
86n0wPGdv6h1usBOc3qKNn0II2R3BlYaDnzmpb+qLXenIdO7TjcaXEjJSB8uP0/7Akhj3pPDR6Pz
6D/kZEhdioTXa+qQn2W/igsq2cVlP2JlXFObkBGLcNYGrht9PgIVI353fl4xco3a8SvPTnHnGGBx
R4q+V59APKKZ18udHAB26iJi9OxYsSli+SuPQRV8+YRs4lPEgNT1kq7spIQrzbxBa5Y9YWOr3IXD
Lm4T1m6+XcmE2gyy6tsoUgIg+I5zvLWKt1/ZtES8VW5pn/H9tO8Qj5Hc7GPaZkexmZBxrMukgwD2
Cn5j0sP0ncgg2MAlSOGEGArwKl2diJCdw8FDRCW39g8+/FtG5wYafc6LSB/iWqMpBbrwKfOQ3c+j
jCoGcKuKsVNIfhF8H64ZQnN60rmBjNYzkpD0U08QOcf4JuBhR//wbLy4VYu5dvzbnVBB/7nXsqgX
/st7LhHDWfszB9MySiL8ZoCUoZgSuXP9eazFECzfTLrch4WD+PD3E4zq4T+hIJtrY4DkZ94xPa/U
iLLiwDNAbdXXIQntrgdzv8WKHj6zDlyTcMJRV1e01MBCOQHCgUYV71WBhtPCnZmTSoLrbbCBHFn/
wrcOTrxnppBbL+kVuWlEIXMo2B7H5rVYtdUVlwYsVhHADKlYcIIbchkTkPdqzMniLsQun2YQC2kd
S/N+YhAJ6Cpd3WRDVulqIjddhPBs2oBLJp8or+a79VUsw6b764KJvaazsLQ/nCo99ba+omwXm2Eq
YH59IQ5lKdiGrnChJW76EAvM78pNdSsoKm5+fb4MqYYipEN8pOejKqR92cL21UcVGvAaQBuVpOZF
mb7oeood7JwRGR9JWyWOmtMgDaVkl97+sLYU37OukTVrjurvp1i6PusV6u7PUf1Pv17oiYbQ3ebn
Vjtk1k0bEbdeyCxyLF1tpZIqiRjuyryMy6slgnmQTvpkImoidjDNv8dmAHZSn7LZulZTAlcW8Ysc
k0b0aGAmOPR8azNFuXrLMc0F/95YiZCgIklVPT55VZkDctHyrhTLOZ63+edlx38DHn0jIKeZxvPt
6vhxxETcXVLXi3UZD3L82aU5Iq0+o4C3UlKn/O5dvpCO4+k76MhP/AcYHQDgk3qYQM4TsQ0naaY9
Fz0nV7iV5FMyLK+Oi2IGxvJDWDurAQcib8IRn8cRDw0pTcZ9GQbWzk7zzjQU9zUpWhhgFLOnuL3g
kcD/+JEqQuEtdciZbp9wjN9OatRK5RRxQhvJQRmA7naJyxMDBhkJ6A6IhcXFokyy5u00siHOw1LE
/nN1XVgyRem6q+QrW37JftuZ9K5bbddzifV5kSrHC34mV+6hm+4PGkLz/I7GUxhSCkm0Vg4QC1Hb
hCU5am9T5X7TqqbKWYnnVzyzte5xFSxtowwWCFaTW4HyCCHeGjGkoDcR3vOR1IS69QciEi2Vxs83
YzxtC064dg/cs7fSO8raNdBeA5q+QZNcrFcSXPPJq+CZMbKqdczx0Z39Fw9tyAYKxMPStsfNq+nj
yOITp1356B2E592hlnDTrSQQH9Savr1/QpXfF7y9eD95M6nGbFd1kaYAnJzw4ngWRZi2d6ULTrjy
P/rzHtl0Ho+DlRM5Q9b3a7SBUaF0vZ0FLOC+AfS+BZwA0ssKGvVW8cgFDArjILkKeO+TzP1zh732
KJX+BQR9RFvtbrjbTjSAc4NSenCAPlKUtEtjinDZHo4XeXlRx5hM6E8CpFIx+z9EKlTDFLxUL5wY
EU4+ANF5A0S2pMBsjqjdrPIyyfCGKTFiZSW5RZW8hehYi8G1hEzzfgJKTGvBaHpIKSW+Ik/QPiD6
3ZNHztlGJWzAkc/pe0reuPoaxA8zUIrPgnfdmdmWztcr9HtRj0w0IYT0uiirGtkrIxozkN3jPXKc
/3i3wfYjFk8GnRZnp1kewN6jjFe1FGrQYHLHRXhw3C+iO3+7MibNDI6M4DyVbGFj9q+m3gqqSX3k
GtwPzi8luEu7LV6/Qkr/UqueOGd+Ap5DQFlGAWQiwhWXkelEobdO2q1OoaSObE4B0RtdHTXzNsgw
KC70A2T1FzgL61uIoFBSG9FDKCzcqCa3GuYWAJDKoxoTFIabBsiIaOk21xdqHPd8V9ZmO47ywvfI
f94Eq7FcuwJAyx7NoWqimKKtE+AqyQH7rLD2LTaj6Dt1uC4UUi9dbjXdn37w0n2r73IvZpiYde5p
nha+toUp8IWR0vRoqIgp3yyXLtYm2VENFRJJYUbRHWIOOmyhR7JT8X/6pLT4+jrylVTsG45/N7K2
DzlSs+Zl1QZW6CGNRh0tIs4aEhq+KKYWT9Dgd/bv1hBBlmcPq6RRk0DKQy0/SQIL03Y1uzagIoln
mbhq2C0KfQjaXDxNRVId0W1JxWaszQT1gusf9PoH0sfaUSMfFLkhDrmOTza7tCe7KYzhN9BxTlki
tFnd4zBcaC7Zg1nKWJNA+Gx2Jxz4AodQzGXdZhr+7KVJgyEYH8ap3KmqVAxZJupnUtiBelkARTGO
Cc0ICA2L51RP37uERbQQ59G1ps3bMcdWac9k7krObt4XPjOjul0EkL0Tng2TBLj9ASq78fG4GWji
o9bVYuoQVb9ua5QawEZD7cXXUeNjU+/yGGgLUyzlpKDrSJ0W3VQX9+FWKWpcSi1RKyk4Zu4y+24y
cNb2kPoBnXlZe+KAe5Ckny15MGLSdDBRRVH0BIU7vm/hHAMBrm9Fg+yoxohBb7HzCI0I/amxUTlq
YrU0xFcD4idGLzVtyI8es4K55XCitdMdkW2lhdNH+N/Et1Bq4K6wgXgqvoVkH0e6GHXYKw+1mu74
fW55Zuqp2I94HXPUkQl8nu7mRAoVFtVgKMbNAeEpR49oRARUhPwkXqdGHdeukfujPJcrR1w3utah
pTaXRBjsKttLxiplVwXgNxTT3p40tKg1JQV7hXSAyhKfM2Weic+z5AADer4Oyo2/GDN89ixFoGoB
3EeAPDW5aJaIstzHFZwFEBda7vIvZ8mXdPVdmuHW5oJjrcCgktyozqJ8LqHMgxZqXN8+BIFvZvgr
9MiuQKe1N5+RvJDPIRVRfQKqYvIzDVYMbhLbdqBiRpu5R2vMBiM510E8zRAwMgaFzCj+GLqYTWXS
tIN+rKaSMr+7T4i/40ZX7gEJJXK6wd3C2S32Nlc2gyNAY/6JOw9w4wRuJivwyM/NWR/qNRlY0wwl
lPhHQ4+dxhTrQGu0rE2/RAhCqHyhPQVjHHkZD2bVjUobHJySj+9zuybiYSOqd02VY6bw+e/Jc3x1
MzIbjY3DJsJovhrqUKsrlBvJEfen+H58A55pXRmyQyYYLHY8lv6nnhEbhbOShTG8SleQawdxg41Z
RODQPXsASu64EL3xYEJc5hPJTQ9X/Vfc/RsPJaZXTyxDQfOl2SK/wJ4xz7GigXqGrQydzVWWtbHX
WWW3fpbxL4RPkuBaqIOJjYwMWi9hZ53bVyMIgJ2tQg0CXSXVTdHmpMGUyygej0P5rRu9s5aDvC+J
Wm+yKSWyF523KIM2P7eJWTdX0R18sAlHHl8SxoU9jw5u30fbbGy4Sp4yCN6DXqLuXc4K2ckp0YO4
9kbTEwOof2mIo9/Vcd0CkNClEfsM+RoH70h2eLCh/bZXcBp0WZpacJmmKoD6HQrXrSqwfKYU2kr9
WOcNp+7VN4Wjf38wevBVmJMN0YMdetcFrcR+OduC2of9sV/gkxuXSCY7FGFUjDP7nQ/mOnETsAGf
mTRiPQ2xz8It69adMPhBxG/SQ3WRUuRgRAB6NDa22d5J1twGh7Of6NHI/39OWbEWDTHQ/7bx/vVB
9i+0Eaopx6k53yyO2r/JNwGbuat4F4/6/lQ1KFpn1nvyL5l1QhV0w0XV6Nxq+V26NPUJ7QQwKCl4
g5j/Qgkxp5k1NPs4p7+ewsSJuuDKwxX+kniRSwSOCTuPsnr8bgp08vbKmv4hl8G+m0uqq3bDKI9w
+FZ4pp4GVO170GNv6o5eQfsdVFmCgcpNSFQGUXRybRScOJXneJzSzf6dzbcFuzv+imq5kus8qH/8
kY/fXNFGgw6lYFSkQ03tYYVRFKmRX18o+qgtW+x2YnPqGV/tWF9WxG1yUVf4qB2jZg/8jX8lGedI
cbaCflNalhBR9tv9uQjI6qe6I/FiYekKUZVDg6QCO0/2gU6tz/bayoVVKUzJ6i9XAY53vY+fyXA0
+pILDzrvcD2hKmJucVz7IGUNDlJuRJkNE1Iug8L9R/TdLTgkB0HXGlaYPrJrB3Lpc1wCo9jS9XbT
4pEbzzfX46iIaxXhPpNHQX68vWfdXhE3rlPQzQSIIkW5tOUNFLXTqmiy1lQVIllXyfhZXGeRS/k6
eBJpPiGAEuZh+lK/XvINKfPjTZTKywpZ4Azq0hu30mJnVlZk90qsyL4l5grzEf6A3USr+kDJGJss
PMPZNvu1/HCA325D9JaeoG+2VsRMLeBc++NkE8AKuf3jcluvvehfnFcupCGqHSBJZcFyZ8BRKxEe
K1TH6MwxXNxpkSoew6M6RD/aT/4wxWX9JfwuMHXUcIWXDbH8AFIQE8VFAonXXnKlDnd+MIqmUoRS
Y1++LN/VZ7bdJRC3f4HFiY0zgrk33/KWdW7tVaIt0QMpC+uOYj8FfgQaPWdCbi1njXYsfBrKZtIQ
42fEbLh4Mlkv+65LMrW4DCkhhFV7xm4uNe2tlymrT3iQUPlP5lvwcOBtxcTC6bZqhsZazoB8Zwnr
r4bIXBBng/s43O46E0/cWvHqWfDQBsb+SiVRZd0arS5fOCzy6hZM3Js2TRI62h88mDWzvuv/KCBu
PnhwbnmUX3BVnn/lSUpltNud0jQ39vea/TGrhQjyKCZsNb34RNixCcyFYq32/bystJxVQOqDyhCo
Vtz/Sk79DPuHs9sEFCyPVhjPVRrHr+SPPitCFNffarjbA4W8f+Cl3SZqcZwQa4Ur8mjdUY5hZL6f
1mJjCN9i0FUpisRh7ZOiCBNbnz83ITX31zmx9maKxwa+uue5Jugp27vEcE87uudU64+2Syawf5y2
9ks5u67+sHzDARUF7/R2fbkLpFUYvmlUW+4hoUyY6+YJ0XhxXixvlOsuEhlh53nHb49p69p00JaN
H4ruSVz2TfKiNwVnuNN0njV4tp2JXTB7U1k7TNVl+2kW9fvlX79wsn0ST71Qhn32dklOgWeezFs7
3KblfUr/iYlCHCy8vAddigIE66H/qmliPdxghiI3fxsa3MnLlUtsksFAMTyegs9ErXX2YNBXnYXS
L0T1cmg2K32cUAbZLRA1oHzMlv34LvNfCSzOANBhil96LOpitGjdF/XUgjebk/HqeDRzINVzcZjj
yRaRvGqrfCzOg8J0JR5UOCzouRcMGHQqLbXBcTTkFShwfm1T1UjBjpZ/hhUyZhlnX30lb2hqoY00
UCRq3R7ft4gDMIZbM1mfOCibHhN/FYlQHho1NmcB6Bc9SRTl2VLR8zkaggFetA0DyK6aK3N404V3
THj8gIZ2xTIQrOQVSDMqy9MePhN/hWW2FrsINzCMZkgHxC63aNCFdVXTvQgVQC2A0/8uj6JuKQWz
kaH+Vh8BpSsWCMUUSjVE8Pqau+W+6dJ4fi3WxMMIq8wkMQPiObIXpQOLaDXkbhSeKzGYLHv2xrdT
hLqYc3cYe/CB1kQ2fXt+f1RIZQLzFY5KbobJN71JhIFXrkpMdr4mlRrViM1YBays+x/Nks8u+e3K
IlEuEZ8Epti1iWILPgPI2b4qpzFOB6NgmqPAoonuIbaX81lpSU0ssLw+2Gd14DAftqvrZ76jRpg0
jkoVJGoITRetXnon4cv9AZ6SkRfbrQ8S1jMeyDVMhC6wVAUjd8lvHsx2mfPc3X37h5Yl9/yyjyCP
1DBP6bWkeovTBSMWdZnLozLFlZuyrabhlbsEWTkJHFDOpSCRUM6eQfcmIwL2dAIGg/oPFWWwIh8W
i4t1OTgqtNFzba7KI8MltatDMbImUE8GGvoUSURu1e8ktgbfgf4/80X9Jat8rg+cCdFyz9YM7ZT2
bRs9G4HkmkGQ4XwBVwqaVvj7H9cBT9Oj4V7GZYWooj+myhVokkBASymeEX3bzWjBUJy2qtMPdVgP
aBnSWzoKft37JRlJ6u/YhCKKRqEtsUov28pOjw2erIJSFEGi9E/tMGU4j1a64TpEZW1V/LZenKuI
9lx9SAK+T+7NgeFqwF+Jb/4ItyBNH8Mcq+KHOhea6oydBbvHiyvz9yCOvcBKSerzl/xkWKY/FNw9
WYa20X23zXIJHlt53HvWoTYFH8ivyWLxxJJDTY8kSPl9oWr0h/lWp3M4CNJUXlyht2ucZ6H+ZhsK
YKGRBzhdNEqHEi5aNLYed8E9bEPQlx5JlNTmA8hdGyULWhRgqopKg2oDUWhevrHbOGQuF5PKoSsb
qkugmnTywNR0BbDCd6IMbN3j2NfFGhlQT2ZMMWEoRWzXX2JTQKAGGWkGfOpzBWXfa82K+l0t7Ng9
qXzMqxZbKzKtuN4g0+Fjf+CI677Jav6lZmxeU60x6pKbO76R00XMbsHIes60pwYZUOc7C45D7cqi
wEALqvj1OcAh2cE4fP0SIQH97qztZ2yDCyUaUakxhkQL6nlksMcKCgPGKCM6IqBIgjqBjQCOH9xl
Qk5f+4mNQiQN//9YzgwgHNucpiIprzOVHNuiK+eJ2eqolwI8EagUQS+4pgLpKhFDo8R8B1m+uuHr
f7oqLTOyxXi3MzAKLOCzwYdjjx222wfylTZmvzSFTHR66nAvoCKkmcrJSKyir5Cr5bX05GLJgu5G
pDvohMb2osmhS22aG1oX9lMUkHIxBL9ZZ23KqM6ztMwl+i/mwarU112kAqgARxtMwp1Era11+e1O
z+BYQyoZUj9wGAHc5sV45fos8BPN7ZEOhfCKYcP/ZMPanHFIg2SUQezFz8O/pvj37V7V3lMoZZ8M
W9GlZXtKpWdvnJT4WYIdKpRNV5vUggZ0awSvtqBncVro2reDo6dWM7Qa9mQyqaESvxIhdkmFSV2s
wkrNrA22w6evpXtqxffXCjHO3YqSQqavi94z2u98BBQXM/ahU1rg27++7GZ5ldb3bpgVnVOkaTD4
9hhL+44RCrFIfq/cypGu5gC/aeNeqhRENuOsLFTbSArkdwKxqGMhx3dqR2ApO+SQJZ9LFWaZDmXy
cTBG7P9nG8C8PzHV46BCGsSiZ6qndR6J5UINdq/czMi76rRsKTrrfsMccjWSBz7Dj0DMAxzpaJTD
PAHTpGXnIVcsd/8QQaI1pAQVObZfDsCK5+J/GR1vvOb9JiznFO3ZfbYUa7UP93qs6XXhfjG9ehFS
gMhozruXJvLH1Xi1s7OyH1jQuYGIzc9ilrm5XjdZ3RWO0YXFqbyi/Qy+15/T7WQTFOeCka57q+PM
LOCHWFo4YfKb3KHbaVsqQJqaSGDbrigVzg0aqTUqXr5rfI/Gmr+epPBlg11KZHWfYdwY9XP2WJCL
4lbAGv65utEDoSd3V8R9VE6YubNgZ8RvwgmYqqP20oqtyxCex2w7j/umUJlAXqr22lckWu4eXx1M
ISvYH9WXPZl+DNZttiLG3Tg2HyhRDDBQfbQ7EW4hF84Rn6Tbrn1uNHNO/vy3nDHVN/MQY5N92uEh
/YFt0D0Ez+0D2h8oAkClnXSKJYJ0iW+LH/VSzFRbSZL6vobmulgi9XKhOq2gOE/FMMAFCUnF1i/Q
1jqh8m0s6cw9Z7x27rgKdW6QZ4xOnCLeYfosiOUUZx9813f9BhzU/KtWG0aYGDeOtxlop8J3zyPS
/K9P/urekzVuiNGiJFGWHyvArPPxEVcMu+Xcc27cGzlhPbhboizS0FPptCgr9esBpXp8JLtQtLsJ
cNcbm+j4Jm2+V/ZU/ykwEWeD/j0IFjjp0vO566cO5e8L0x/LBATAQ4X80h8xBAKrzSKHS1HYg0R6
VhP47DHTRKjhN6GxQPXH/nA1NztFZdnMKjXHeQBfTI0CqVi1I5hj7nu2ZV63QD6EBJZHFH9W8tqo
JhhwTartr7DrfWWswS6SXh367eJK8qmXcf7/V+inbcvQoydWltFrD01mhCXpOUC3HL3CNkhiWXwM
Rn93WsxMXsCkHDIs/ObyfpwOA9pYYmVf0tNP8RUdllHh2YPpRkJfyGHUym6hKQNfdA1aueDIsxmU
i6psbiMees+oiKJFyNXiReR7I6z/3XAIg24ImK3GIQ1O6BZl9fzp4NrlF4MEdWQgEjgWCwH1hsh5
YPRegsomx26WKQScpkARhdcQRtUojXmsELCfHNHEl9kg4tgn4SkQOrn2tBVJqFtufW48ItzmBWjP
E7xC7+RJ21etsGeJ1oXKpGh/HKwdO3O3V+CkLX12lWZAh4zjLwHoDn+V4P+lq8VP9u6t+Arv6jXT
r1WefRCSu5nUbiOR1EdtRw+vX+RkhYxupMprh64PXrotSYNwl/cChLmb2zOOMf/7IGLEuTTGhRZ5
b6O3Ezd2UyH8UVfFHZIeL6N6KU+WWIFjFfHC3neMap2Ut04Tf7hJmq33ufTODqmiudY4WgahvXjH
V5yTF+CEFesCSo2b5YfRrpRKNvhuvtKl+V6R43gWdmZGh66fIDEcKz5IRLvy2tYwIoPZN0twL48q
nyQ8Vtp0CbYk2HYSljWV0mF49pOBgfZvsOFsQOg3IWPP6O0p2efQaRtd3Sq5VYfNBgf3xzGhzO36
JSEmH0FtIlOlDze3Z877yHUE+clASR5YRs6HhBqTSdLjtFRKF/p4X4jtf2YM2W3B5AqZHmDUokZZ
9mxSE9JLsWV3C7zIP3KySPOuhb+NaL/F8/fAbRv9u3LzGGeNP4XcdEoHhC9J4CA2pKe4qVzS7IfO
laA+QuuUxMbcGHHztThHBqnl+D5h4ga+TszCcs062476FfvsauOWJ6K6z/fZ0rDvkKpWcOHTKTFD
0eBDTZ6AR7/AIs7zmQpUyCoCXgeMhcLAJeMeqKaYvISd7sv96/DVhKQ9xWb4dP19yuOu671PPGTB
e1CHUYzIQhmbeWXqCGgg8JOZ8sltXpzUkn6ToLx3pH+B7J3TFifDcn6Jpx1jZGbVwFedZlWOO//f
mcwD9dOdNGXcR8MucJBONDG0Co2c5rMWLttRlxUqfPItV0umiJ9RgUadMgk8eRofckDKFpftIj+4
a0VxMTqyPP2Ql2K+psKufgP8i3+XZ+ZJWfi3C96eqLJxoliVpAEdg1bPyRA7wsCBdOvudIDPDSNx
yDMeeYBKb5rZ8fLAB59P/Utr6o4IboCF0brf0ksgzsefzIDWY1djVvSPg10rlZuDZ3BoYgBWCtH1
P0dJ/b+moNKMC8NE6SXxKV/gNxZcJP1koifIN0Q81AZ6vNDrLYV7Lr6QDfUOhjZqNkFwST/5z3Mt
l4NFVcNeDd763moq59M96VcREYr9uYKrvwCMivP6Xd1lvMnDVMBV73dwa91uID8QFbBVd7wPTiUe
H6r9m813aF78lds9L0lDSVOHNxxvRc4nxhcUaJwR0plUiYK9oEICL1yOfc8B2z9f4bONnoNr+a8o
eOf3afpr3yKO3ogJNllrK6f3E9CPDNpH7J1oSSDEXjQeo2nBtJqLUgCKQs8cSB77dPEk5/SXqKNd
JAyG8VVjoSYMeXadUwrq7+H8FFI4oz81YqhYLmJXQGqYYrWvX6hVu009BYUz2ZVbRMbQCiOsQYx5
MgByzWZ/vRoLZ2hrA1mV+4+PaieTwSAyraPiBoHs2iLtC5VnnDxjGeWJBmcKT82e9oeU4q5rRVLG
LO946ifm98FZllJ0OQmcrv3E7RZ/CzESOc8pgGLo881t4DFrP7Pfri6NhduoWjDKUhlDuvy9pi9r
rtJLuWKD5Mb8R9Qrk4TmuFMUDkLtCYGVbsOyMScI4TZMXrW+sCeZDCkFy8xBmdub9zprZzupx3uS
N7mfk7dymg6m1Mpb0DMmrZM/D7oTxrRlU0+2mzrCJ2bvZTPbBSqUFWEDnVXZerX5itdwZuB+41H9
nlsDVNd7NWc54JBXC7xntHuuvn0Vm1m3TWGWbNe344MvAH53t5bmFsYx3hKmObAREvXchiroBs19
62Q0DNu4Eao1q+VRQDphbpTIIMDSxixa91egw1xrYbby/NpAb0UgkTFhRPLi0A51s3Riu4ohdaIS
hc2jQ0pdAkUVkH+ghZLvMvZ4IsRajrlC1ruIhl9RZy88+6akVU7FCuJSCBfU25Qv5QFc6+i6R5Kn
nk+HSWzaHpMWWvPzYzmEzOxDAAYceMDbk252jOrRYksc5llOAZQO5hmHWHfpRz05nlAA2HD6uUrz
k8nMxI/8VwdSoopTkAAyhnWWEynry7hqqKuUOTbUEZOm72UmD3xIWH+mXi6jGnxwmsQKqI+hhl/m
npFqBcXlXMaHxAcDLZKwg7A6eIXIW+HeWhRJYvqu75ql1OF6SA0syp1QCxVVWaJjZ2H0tL5WRYou
RRDsSPS2ZC/eY9fR8vMCaM3iTpEy/PcPu4Ujq1tSruxU4f3gp4vriid+7i1Du+lqcTO0IwcA8cfR
Z2RzVR7/lJY6abL+/ypkzBr3Jz1MFBo901uBHNLhoncyucVcPhidLl/0lcE8eye0QDEoljw0w+DE
+G0HGTs9d7SJhufZ1s6yOy6CQ8R7hLzugrm5LU0Bk181BriHuFScusIBPMXilrN0ZpLz6nUhq96c
238wnS7WwtAQ4sO8wsnmmAJf7RcfWXIumUG4HEhiJTHA33YbXDalX2qoXcb0et2TqV7Bju4r05UC
kL1Nw3hMIBmCG1mzQqK1JFc7O3P8jZnTM6AjS+sNSdYavkMs4MlqODQCKUNmJbBy3hUxpsoQ8iCy
bp5HqxCPSRD/MZCHpYZeoO0IimvhLmefvAQlxqedvtE2MHGnLdCj0IOtDSKSF5j9XvN5ykun7WJo
ysEmZRyFMPN9BcFd7qRRZ7uO53QPEXrBuaOi2m6kUJEL/cGE82U5nJD3sAsOXMVnm+rpF6q5u//l
lxbp+MXU6uDUhUrbrKDwjwhJpc67rBOsFri4ELV+7g42t/ndHpgmOd8QTJO3B9dNjDe0Z8uw5VQb
O5F8kkxeluoSXNKPuwEQPPc/fsaNu7Z0BhIDkF+RjxQqPXCRz+/bppdjMVYvrVa3DVFESO1Gzo2n
/WBmAbzGRRkYFRGDoWFkepGW58P33ZiThMzZtG1KizAK1wgfOny/jNNIlrL1mHmnarwiXReDbKIP
551vJQLqMuf9rD2SuLx/hVO0WSnEslb9r7LYXweX0zmjQA2l5+rGdBnFWqqFWjYQu38OeW22CElW
pS5Sma59vyWqXtlO7yhsj/DShkw0Oo3OBgOABHy40f+rbPrX69llpgHZ3nfbN4JTJRzspjbvvSJV
citFo8dDPghf75p+Fyw3xF4UNo3U/IZjXTdFTTAmozDjCyOLYHJABazOkoHTMABLB8vYilNDJrId
vPLigQnWkhfex8w0m9bKL96/ISA5r/DowYH2u7zHsfb9CW9YOOmxkpnQLox7A51Cl2EzDCp4F/4K
VzewEBkPWtw2xTvVzsVvmQXwp+jgGaaLLT1vBcfw5AxPHfBydvLhQVQADACocLlAAHrO+GXpQcdQ
ZapqTiYMMrEOxQFMUnLjleSToKqOFjyoikeRHA4ZIxxv7Bdby1nfG96f9W3f/zbcrZjuisXgAMHC
09FHHmCydhNrC/9YINXGSY+X8wl58QfGqYuTC/wmP73X8gEBp4cwoD70z9ONhLiQA11n5vNFNRlF
FsfAZYDkcQJSsmd8Ke/gAfSaaODurw/AeEiNPrAzSI8EiX8lUZI3DrzVaNoKQQv9sORpXAEg+C6X
ovx9W7/hlHBNFbkwxobRQR6zfVTeo8u2qQc1DC2gaZCcESzbKpdDnWqMfqTrRqQjcl5wiiVv5kXw
4q3CtN3mUWrRVuWlEehZXyMJwWc/laDb6Pd3SRhv6FevDDOExQfqsOzhWn5sfwpofmZSf7Pn8KiW
RZ0NbzjfsqWEimwsK28A3fPo+1VtL/FRoHz90TRUI3AiamQtRwk3tQ0jewrqWUHUBvK3/C0w4Nk7
1vqBMj79WumwrvBT8B6BJMhCeZ4ukJAIaA2d28sU04nOh1EQMIWZ1WOZloAA9UDCGLfvG0cdYNtK
heuC4RbkM9yPPYFxIjx0RAj9HECrddKmCU6YyGKTSTfZYMDI/1fRlE4RH4NGlMOfCgb8+TfrM5Mx
DdMFNUj7D0ManaoZHj2nNcOYE5niLYNjk/dB1Uvmh+Br+FE0q5QYz1smJDNjhl6u0uwnq0qIrPiL
HvNt92LAI9uOwJDcROMD6Yh6EKLYmfYjh2A+MDg+sDysrlLVv/PQEDfs2mK18+5wiQTZlJXBkB4x
QCcZugXCLWkZffCsdzvTMWLgmJnc5Kgz8GYXPTJqANn3OEt1NsYylanfdfMzczegfBK6X/J/zqhz
nAqWlArZNKIdeuCPozfDGi1skMCDsZRnbqAk3AOBUhEx560hVt0RFbPoQcSVphCoJfuTrhiPxZ59
YM7zrPDYVeFSG2Sz67FA09ahLdQSYdTl+qOZRjpyer0+a6kFzHpSWKC/AGCRZ/PSvZDYfixULQ4R
qnqhJQAkGbberBTerIC6vTHFxl5B3Jtyq3JwVJC/6Klxu/M6TKPDHD9TI7KDKrrQiFZ6dkusEG7x
/XW1u7qRNlLtCVJK3e0WKKoGMQnD4354tt3w9b6/+zO30CAhDvy7uETEVnlFjMsJ4CgH36MwJOmf
Zww38hpq9xPx57i+0da3Rs/5LGnUsdFGX0GRKVuRDlUcZLfPBl2CBKGrkJSB1HL3fuNQLNpHSHhb
5MRm7Ew9ayLVozzGiTb2BIdruo/CyANTheEi4BLV1oe1+P+UW8KH51C7aYSd3kBtFxmJTTEIoXG7
9tRyAFcGEcNGGhDP2WJVz+syvx2cxem1senIsKqmGwob/dkPr3aWYNN/mXgIiDgMlsyKkATjUkQU
nr9aMQE7u9bGzlIm0IiA5Zu5TYXt/2EziRzkpcuJZA+xOIvsMRC92rxoxDJQfdb14iTM4Fu7E/oS
hFqCULxsDfx2k5sL+T9KTSmrUWR3A7/BmgCxvClQLwKFlEKSfPi83A52CwPolL4JxOTe8ish45kp
o70s7hH1ReVTHz4FWU9ufN5+bD7jQ+vPtJxO79BYsLV2QuyKlN1gfRpHg8GtPYQKFSAXEGwTWlBL
fg7jlv8wTJs7QmT6WV3z7hf+1gkVVojwWcP3iNDAzvjNdBeO9xlnxdlpzaAbiBPGt9bsfDuURVq+
wbaJ+KaAwao9UjV4HlxyBSWfkuD6PMWM3obbd3gKzKmk0sKCBnfymWHmhIy8l340VxTCqbtBIN68
ysZQD39i8wzbZYXvxTP5BZVfNwi688+BISCGtij3ACe5Z2bZVwQFyBRKuvPwQt7jNaWesjIwObNS
vd4Vz/LAItD/KRBm62FlDwyCBUQnfZe3MKn89cPm1ZURc2qBxQeKDEp98Z2bQhjh3QTKkK+iYy+M
vJM7zHa5kefUcctsuaCZ6qoZKtqd176E3APm8X44C/vYArBODX10JS+fLUUP0QnFuHEwlyrteU/K
0FKtekh85nQI6Yh+UILshCCHK3ya+Fnb9c4nMhLoj9/PA0dwtFCgcigRBued7gm1GE/uKK7AbJev
IEbjg8UzT3TB/2/VfzBUkzy0R8x2GMHcTCR6PcsSGEofeTqFjFq2F25AtN7xHN3RRGycrVSFlTSS
HYCGoaOnP876ENpeHE5PceGHrLSTFWoxlzpeYeu4d4GjPVYO/E94r94JX0llB2K/eUtzch9xZPxQ
6VLPHOjhzBYGRa2jcYbIjn/AzUpsrsVWIdUrAWfT4ZPDgRWP86QailOqInrNQjtYRFYGCQBgcqQQ
IZ3l5uYQxWa90208vLEnYOkp8f3TO9PU878lLMk08MoDmdMArL8aCWxwckRGhjk+zm8aB13fPOaE
jhmzzyF8CNebz/hTFV5hXXpnjhu7HQHFZLpAjljYAsHdyHNc/L+pHICFslTPZJ9xq5v8kWuCF9hU
G5A1AoQVmmOo45N5FOWvVhUC1zGSKjIuEqBkQwy29cFobYp/nIrmkbICORJaOTPmnz9rkoDuJWgy
HKRdOXZYW5Z6jVuRMHSB1LjJnGkwEFXRpUiit3i3QLzqP/4jlH4WYBAdqfIYuBYjcHA+YX7kL3jI
wf/ThVsH4jWKR/HCmo3NlpBnZIb25sGoSs+Oxy+WId9QqUMMONeGVZCs4MHU0nJpZyqB4OmHe00S
Dr/9YW8kRFroROI/gmk204/daxToag2hwah1sHSguUiA7TlLmVvwr4I9U2PCnm76J8D01Ar1WT11
CSzdyhAat3bOst+sH420he+gXReXHOAdKlPUZDKYQBtLaFJ8D/e9mA13swyXc98imkeIhYwqxZIY
gwjfWkeF15uYboePorGwow094XU0WZT9OdihwXDmhEzvbbBp7gZ3OxjMfkzIEqGxYzk/VuzlkJN3
7PoEo/NtM1j93EweChqWrwDOWNT9AAzE7jSGcKanvcWbg8sinBxvM+PvpFgJ6cHyaWZ0TVazR4nm
Sa7W8A3M3u41p1SJVHQfk3vLr7w1zg0NOfGVpJTuxBgxXMfZcRv4XhZS53TlQKtCt+7CCdQF2qQ8
uQpsq+rWYKEyBAvQesL7rDHd4amwsLxos8PMJHKm3ixJ0P1fZbUKpnipSPSUGWMbapX6Dv0SZTZt
+fYOIpaW5rhJ1fFEMFGFqN1qdP6rabzhTzI7BMpcRNx5QYBoJi0coB9pjNi2URvoo+lnWLyZUNYR
j3K28Zfp1q97ytrqeXCEmBLH1PdVAEmaFrV0qhJCyUYWVPyGwYTtooNGnaM5iAf3Bt7t16zJuK7d
C9igEKIdEzqiKt6NPfHkPlZ0zh/CtPGsjq2YJSX4WTC1He+0SwH17gKo74Y1fkIqjWlVmHd9dYOw
hSScCo6kFlpJjQyWw/g+4GjWtmKHJwNfJ8mvAfDOSewa5QOy4B9HGg6QjHubgAZP820MBYcEQPHX
7wYpNXv8HiY0NcOime7Ag333yb3FCzzhK2P36tvN/VDX3sB4gtPwRcpJbncIFP9kXnnGfN0407kG
Yyw9fySETIWF3X7g0xVLzvWsnOg2kx1I8b/C1abb1tvInVBNsbUBdD183SrfLqLncphUrHndQU9k
4aDqhWVeZ1dfl8AdXkj9d15FXC9z+uov7Tz6V8IK7dplu8Q95v8xL6eZZhvvpctjQiqhIF3gE0/i
Uao2M1UvOaOjUBTVCev0j5ltNSJj13d1BC3ct7Cr6XeyYKr0CYpM9NzZSMFJkE8S2pyfoge2GrpC
7FKMCeZWgVXuln7Nz0iBvtjio2TtwTeG477f4l3oxnXIrcIWlWu7ERaLs/br1W0vJ5qUJRGry/ij
kC8AZKfz1FDEyrW72gWaBw5DnbVd/ULwJ+DK8gRPDYHZ1dB5dGrAgtvylV+YbDFxQhGLiD+ISH53
jtzuA0PLG4W8pHNsn9WCZfj5kdARwASmWJd1E2bt5oHJmJ4EVUPmCuTzAy6nLfvsQNozqJtFMm+M
cWFISfGhltEus0Ssk2PHujYhWt2tR3VCs6g4HHsO1jsu5BL3mhasm4nLlqtbRXinHfPOo4pNuK/0
nsGlZLuq+XJ3IrfXHQfXCFqtKXjkW3dR8dIe5twu9SBnFf0seux5rEMeMuXDga0JSfnVhRQgqjdg
0MvF/696PUM5cydmQv6qnzOxq0KrMxkNEaWcKRAE0wS+Ocp+qbcQY2EmWc8ILP3DPkorItx+nv0/
uhVmNm7bSTxppnxQUmp+noUtlhbBFrQ9Tm0gwyK3GinrO3JTUUNt+rmSLckhqJYtBG4qwo3FqrB7
X824rP1ZBzta6rguQj/xFywL5oD97HYgGQ0rfBBDZEfQeXbHWQYgA9KL6pb49gcYKKlD67kIepbu
gL/bdyxXahWohW06Ol13BPINa5ln7Dv2wCrAHO8XConG2YmavAi1QsP3uy4bjdWfIYiavnbtxoac
FD57/Tprv07zPRr5Txo93xZAd2jdvAUQsfryNak2OFRcXyOK5tGpQdQe3bIu/+r0iytFJlIVt67v
A00AgwQ6FKXkIC7KUY59FaBlTNGa38ofdIqr7FSVPAY2h8FQhKDwYOeG5DXGNFeSWcUCk4WS/Zh5
wQ1Af6dvUqVhgUWYC/gyb9ybuzfRBIyhlUyovtLG9Av0y2ebggL8ekFq/Ilh5k5OY31MM4Zy7c0O
iQDb3gd1Dpj0WTe/DHEOVPj/TNOcerNazkIxBTOVN8/FOmMP59WDovduxHmf7FAtgXapZUdLz+mJ
zGWy2etaeUoZN3YqtT7ZqbwIcoKMzy8Bjlq4AkpO/T3/FXwq4Yqbm+/jnVyxcRuVUkin1Us9FPCO
OnS8uxIBhs3LTZ5RVbpAtVKmywMKl9p3WVP38yHIFg2yt7mOSTpbo2FiUZh0JZgmwmDFgkCbjqyV
wK7vu4aAJ0SjibKDUuP8SJKGXDkCIsGAV+ESOoVACYfsMqQPbeFDUhS7b0ShC2nYXOennBZBOYkh
13iKZOxpyTlHf6qZ01a0T6/UZHEi7SKeqlu4LfLxzqbO/Wlq9VyU8bFvANo2CjghrgvvphdumiX4
S1bsTaowS4GU6RREYltZdBRFhi3d9Vd5iEH04xgnSewz2sXM7puIhMxT7tpBTtGDqYcByDjNxDKX
FhOCo07B5/zMzdFRPRuqFU28sFlwYs8ik08wGHTobSsH7exTd3sl9eyNltRCMZ3IxU8R4+LzOfAN
Ao8ehNpIXm3mWiwpmAp7zn0py5/3k34TXy6CYAsRkxzCwjcU31T++7lCxUla0ehmdYW/N2PDj7vK
X4ixObg3+0xXdV5oFHlPSruh04srGAz9omrK3mPk7qK0FPlB9x2LtC1KiKvXCpR9WagmZPpbwyV5
waqFPkRD45Y+wJCe7y365diNzLeEIQIVdzQbXLjIp/ShboLhtyvEfm0ymk+7rWEQ92Fpf67Gr+69
cGmrOOimhdm7RfgauqcyOJFHHmX2vzzmQILiJQOTaxr4/X7h3XoQd4432LsfHwi59VPrAcmt0VAS
CkRmdn9D+IUc/L/taNBAZy/Fwbl3k/VDEIrsejUwNTaJj7khahmBjQ2adiAmvSBvJTd7HrN+ckMs
cZQ2u1nHzKEvjXmOzMJ5RsO/2TdioxuunBprRj/pAdwxX2YMsQd6MXy7EDI8yKhorJffT9xzlwSU
tl0HaHUsxDLw4TbNm68b27rAoYeBbkNr08Ih4M1jmf7N61neHmGyjO7f9kW1uNDKRn7b9//3X9u+
3z8VZ72qL5yt4xsLHQr7KLlMpeRbDsgSAw8bjiB+eRoTY89n+D4koJ9VpTmeeIDjFIAlkOMRE7lb
KXs9Mzg3QJXEFo/HuQ8njzna38nh1Q5XgHIoYM0DU/nPhOA4y7xYdpCUPfDG9dBpWzzDVcjCr1tj
qMfySKQQ98XWvrBo1/1ThDb8/gF97km59Vr69PuLWF8hKYDPe3HZQQ/mXJ56CZvj+4JIezy5sacT
XLsoV1nR9EVmop7ldcwGXMJDDu4zEMVkFixXyQBimc6p6UTvxtLgwu6h/IlKn9Py9SBI1XxQLL7r
L330A7gVmz3ICzB7x/i4oSlCvhu9eRwn3MvkWAm4OgW/Wuez06zYTeeyOO578vFEGSxhXbTUq4uF
pvQj8px0WWt4Kcs/iv38bCjpBjArCEEGglqYdSjKUKWH+ZuN1+yJJ01dVrcBZ76aFiUccLMSQsd7
hzp5GzXnriQeN+cj1im+ylLsieFhSuI1xt/qUwd4Qem15ChxvTzboxT2hzekSzUrnfeMde9FJV16
4DMHE4Tu4GtUjuq4IC/EoqgklF53g3FE5X6gxsXPQelknkxaIDKDSg3xRXNYi+2G/ayiEGrCQ47v
cwRg1Nbf28sqhkSvSdxCEWFnoPJEfeUWVLrx+P9LszmwHHJOCvP3dYOxyN+WbQUwegkl7MrpQe6d
zQQNhDDuxYI90EqZebO4227yguKxA2QdZCNzYf2/EvwP6ybWDnK6tTPrOg6x/GtXOrz9VQEJbGaS
3Pu1eqVO+zN44B+SikSGrBcn8jLShkG4GkHyia1hbdu1OQnxBAP335XnD6T5IHeA4LgVmNHFzYal
ZQR7urFXGMnLFvJ+/u/AghiNi7jD76PCtOfYOTi+MpnW05N+ichfB1I7D3DGZ0Rsu5ZzLHP9bwTc
QGvQq8DCVjxK65JV1eSR5yWeCXASrVScIK0/IpAqv4O7DMrme7AjRKY6fh4n3Qb6YTcdPRaf2rGY
fPCaRZJD8w9zq3RCQAp2TRjupJWQZ2lxzaT+k9jUAGTcoINec/csuzQitei++sXvrasD0MuxDYoV
5r7KB0ugcIcq0XZYgf/R2Mm2M5sPlAqsCZ3dt3MvenqUFtcDlMDpg19pLcJbXMNi8HrmSLwn1Cjh
+PwGz0f3fbL7pxMyJ5lZHADy6275O4qLofKPCR37cStBhRI4Q6ggoVL0gCFLIkI3dwu66byKYDVZ
aN1b5uHDqEQHf0G7LJPUkQ5NfIAw/+A1dPyZhy8D9nS1Jt6ilYMH1pLkZwlE5IGQ1O3iXT3iSpiX
6kQ8xbq6xsenwBnMUJLmwgP8ctC3MleQf+ZEQOVmXPGRHJ5q7kStFgf6mM2rCDw5nlLw728Cm5/H
sNijOlYIkZP2qa2lh2ERvgpwm/EHWNtMxirBKmODiCIcouaBJGuPKYvSp5cxTk0fyR11N+MAWGWw
vgXZpnnAEPDnYMcyM5v9EqcNf42Yxd8s63N/iXmNI/NTu/PCwgz9YmEH0FEA9gcssCEIpINSkLXp
JRvwulWcGUk/5Nt8cDLmhcOjyN8bCKN6gB0tMhaRDoYxVONfLeZvGC8casxJBRLHsRHVFf7IfYS0
8EmW35hnjWIuVTqC3vn6Xm/mHjVY4hVZbd6LmyJqKGBWTb/Besc/rhwm4FrrtqVOraNG5j/nCsC4
KqJp+GZ4I70WHUH7Ing+rBbVvlsMjmhCNW3TlnbOQAXpeUS14qWGaVbs6gSrV+2qumuQ7MriGuXJ
BRgYZGodp+UWpoSPSQuv4AFuIgYqaZ/6WFZRWIzhMyN+4Maw9xfiX+HlZ7pLwSfyfcDg6Ms56la6
g3YU5CPbj2z44l004I8390T/hiE/btCePqvHP3JytasDjEYXgCvhnqR0nSSVcD4VTLLIfOu9OKXo
XGiX8A6Sm+EzUKcIU6vRzCtqlzLDQP+W8+6jNTk3bZV/mVmI+xDjHQ08bWzaHqn7Z3OyTrsPmi4f
MrTPrCPwoI5lyQpS/ZzyP/wFJkjQlRtIuuekBOACw3raxBjcsuWaInJuOM28UNbmq45gWPd4lez8
sv3/GYKjoAuCixf9yImGYFtwYRxEoGrjTVMiUz0MNqPMXEsCVMIs59uAmW1uwcmX2GslkZvGMHO9
AqDbYqU0LdA4mKMYjGznalpm21kuwY3Tl+mD4IPNqNMlol+/aLDVfsEK6EEJwCEDVHAXSITTzqFP
ibeva0SwZhTZVobfHx+tWG2OoE8lKlh1hiAhbqwSTF7kPtXMTNgbamNN+O7DNjKmrQTILimv+aDb
Cq4utfEdbtA9QReO6XzJ3CFx7mRAAIOKq7n6+hqEnS8vH1IHGiQp41586S8zMFmU1edWj6TTMc5d
APD/SPuNJ/fe7WKvXrXcXKk/byTA/EEME31KdKEuLR3YpO0erAUIq7Ao1GnkUnx/nUTt29pIvQBr
25655uNUxIvZKLLFvt3bd2eU/sko9T56HfUuIToM0+ECtdVkTF264pCZutI56LMUo2VVsJQhEedm
y15tfWrMSacOUuA+4zmwHH/8QRGZw/rWKZY3OiDgNX1QAmlRsaeZLJ7z8fuv3sJpgkWTPTHMdzQX
MZSat0HNbRb9pvMZInozP7ldvqCtCUcvnbFeJAXWof8UXV467GvBCdFN6417jBtSXpU98qIpe+01
Qu+lBowSRdgQ379TzAHwfefljS9YnBeHBOsSsILW3VrBepwkoyARgSH3evng0PTGOumNcU4cGbLf
TdNfd9K09o+4AZQ7ABO8ZbXxNsWHEI5C8qWB57iEZZ4IUGvtiK3+zo3i8JdlPa1InilCUYZHJE+b
uXDCoxykQC9U7q9G/LddoIGyzsggJhZloy0yA1rqBuKhWH3WljNr3EruK5c0PetMphggB6RATIXO
1xLqpGWqv9bwR6DSLp+AyNcWrPCoE0ML8RSoqGEyclx+5dnbJOakK7YgeUEywYgwLX8J/FchhzYM
7EGkZ6eexQeOKsiSDiy8O6Ppx/D0IveRSgccPIOpLbuSznw48AKL2/+sZM4+DDCafPOTM8kNZDRv
6OWPRc3UzlcMI5CtKTMdrixsdWw3YATy9ofUZrk0LWRWMPiNteSZhmKo/6sA2/9vfti79z/baYZT
9S2/5pZsL09lk7h+CIwtK/CoUnHPaLdkLDjCn9pUS+vbghHIKSzNWcSlBqlP0rMkIqdRnbV6W1ak
W/Oe0D9cxGiSfFD/ixMPTx0no5lsmMXy1ZU2JoJFn4ksaEkQn0QAjEdRnCFbZ1R0oSoEdW8lKXPe
qmA0MvYLcpre6BK4AgWzodKsK2bILxKraJso5LaCX/oL6yru6vmK5aE8FmQWX5rgmsMk/JtBFRAu
pciIGwpHzZwDQ3AP+4aJqrS8QVpTpVRYEPvPxCgCrsdmSb6xU774z3GqTGITfo9EhMkupIMYmWVA
Mi90NXthV7r/RyKhMC2ixgpEGS9ZQOTPjk5M0cMBgX/rTzOoW62NxsHUmZltzdo0OY9X819qmJc5
nBwkH5N7sjH6muhzZ26VJFS04mpVDe5czeT7PAjx5lI87BnHrDd1FgR2EBWLorP88ZI5TBuoD335
LRYTaF2Onm/OD/Z0SQBM7FZY9YW74zW80sa2MplpMuvTwKEwaFdXDX11ouDR1DJxfFxb3ZtmX7Sk
33mhwnXjIbboEfCgmBUM5P+bJRmBpYdHngLI2aV4RDFmjloSKHfEC2vXWMEFup91keujbmnl/IVR
C7W0xhDyOwBFjwXkWhJfXyb6ApMwa6TKfKOHdLcci8VDB2qmByQwcJ1EubSGXjYWxgMk69jgWtT/
tz+mbBULQV2qM6XzBkYlNGL3FTqPn9Iee/1jOGYovTF4qyayNYCnIDCvYjP9vMWEAJiigk/sM7eZ
yuRJJAiY7o+97oUs9Y2SNCnDmzAe7mQFFmPobs1I7IQdD7k0oTqG7JxQlL9xbKgsuEhEqsCm+FCF
kRkSFJg8wmexs5luOCFyLjIKoJmgBjavOTTyGCcX0AWuvPbg5kqn5VL9jKQBBMVZN8WhJK34j+E7
aGtiyd4cgKoWVtCXO0aOnS0uuyM4tk4fVbH96khFUysCvbO7GBVqQB/uNrPVoxNp4SzKTYKzJRL8
iYkhREFZzp69Ci+XxW2TmUhlfsZ8FeTwsN1BhZ+agRUJ4FNoTZtU317xZ0dfLEJJoJS7xJ8PMFIq
nfsUUbjdE8FdCrwN1oH/d9QBReVrTvlIdH9iXUrAWZ8YB2YluIOIF5nCXXebIwz2bl4OS6csvj05
2YGqNkH6JIngPYGw+M2GSuTUsX4HCnE8msq0SVioKbG1YcnvEI4a66bk8MLiULXp2On/wgu/KKgq
K2mP6GPcTDjxPz3fbx0gnePmGxidxw+5Q0kGbCGgW++Ta1q9jywn6PQBibTdcu/zo9LAhZdwqqSf
4wVOu0Un90W2eBrWhJ05ZIAY1Z5jd8w1SGBKhiES6oo9+JtbGOSFCVA25aV8m6GdgO2nhHMr8rUq
lJKY4Yh4fMMEt/Q60n0cC/AJwKpryjRm10JKwebhpsLbHPBQ44Szpc9M+rZsooCzWOz7Uo673Gdv
mqQ1lb/SKYXLKmWGqXYPXfpxs0N2qdXAhfSPG+Ig/AE9vH6qrLpHjNt3hG6Et3/NN5wxeyl++i17
oQBqcFEny4QaP7ppYikfyF0dbSefvIXIAuzWPCsTlJc3Dvr/8o7GzLwGWTNVxZ+iki8GwJnLSNTj
mWXswPxbjPTxXc1AZKi8Kpvt4wlgMswkpZWgFNXJccKWoT8+QtUaW1M1n1Q1vvtWlNVgEafwcPGY
HKqfobxp+dkkv1/JCihb+FByKEyJ6xY9SnXryGdgwNrtEebeJ5hylrzYfQNw0IBqbjj2QIFwRvmx
su0V9SNpGE86wDY1Aq/RsBvECwpjaFOwu+k1Ilym9pKSpM0a2ZGaqs7guFFbtNjay11ZFs17bKI/
mvv3fbsS16rWbcJMe8ff9BCNF6TvGACsSYmuZ7zgSfiIk4q5TAt1P6nCYHCtGKgq2EH3M5MHg7+6
+baeXdQkbf7aFcNBrZL3b24MITb3IMbzrUm6HIrBXx3c5KKy9nkClp+j6FOS+GUnkFHw73TH7yXd
tb1ol7psUtQYTbzA3PkPGJSsYeXw5eDnpOmL7fA2PF+QE9h4KH6gO2qnKkqFZNjbFd9oMdOY0ajM
65n1o6aB4A3LGqmFSu+tu4FuM7KgY7cUI1z5hv6oQiaEJcdcBdW1lf9i2Ge662C12IP83rK5kvAl
Uu3dn6i4lfbNIYkTX5Ugc+nYSsrIad4CSXnYCVAfvO4QGJJEc0pDaqV+rYYleXSVEYEQKRmZXyo6
gQggpHfjvdmPxQ0V16ziykqDz1so/JDB7kzAEVOHlu1RPQcTyr5CywuvnVoC2fnUBvsnzkXuOuOZ
xkNBz3a4D2oUk9VQdm/+2hoS4cXTqa7HsTvJ0yofY2dP+mX+SqZzf+eZ/8L2YIjNSGEEMn3Q67le
mMoyV7TnS36W3kLQK52ny7UDVbg9N1wM+8gkhwxZwWfqUC6WzVdvQNhrzpGjSeo3GCYOqCh3cKfj
52t+bXmc2gm2epK/WXTUOpHOAWgmsVoclBffPMX03FmWUGkjrLZk5/l/RxMT3/x60oQ+c7/6HK0h
3iia631WIiqUHg23yUqzvmLrSz3SZ+XAT8jhmEmSOpg4RC74aj8VU7ijXYlwNSRj7FMLJD5rcGEi
Ivg1JMxKJUjJakZLXYaWUfCMuNxWyeIy2d7Y15HXTPDrjfQZC5lOFdHBNLrqkJ6aU5Rpu0AUSMMz
dY9kY9deXaKslOKwDFkOj/XrIZlXFcwV1rtZ1IsanshHYCFH2XQitAH+J75irCPH6p8ReuVqBQ5X
hd9MXY5IoU9H8Q00t2TC6R/yitM7DoEH4rlRyVJto2amxGdxX0+e9DFBrvSUqzenDOH6S9OlJG/e
y4F7YfyO5Pk8IIJ2ORQd2ZSJV8FZ8S7fIC7eNfFHuxpx4YD8eYTIVKHnYfzPvS6D+EnASgXVAptL
NMbDcYGv7gr05PYvjEDgu8UviqRJ0ilBDbwEryC4ArO18eOpN/+PgiTIkRj6C+BNfG8T8u/PHMGC
AoF0QtHqyWdzbMGXOPcekHvS0QX/XtdSaMRPnMDCTlYqjnbdCo5r0xvAy+p3Lwhdw1MOSFB17WiQ
JMnyTgMEXHyI4+v6mNFJiKMd2cHAFJ5d1Bfff+nF1bRQtNZjMDjVMs5IAdlfTEn/nymzk9WZvQ1o
hE/LJ8EzGKsZDy0jC2qBeCt61jh9+7/8sW0XXtaXGzlnBkrJoyyBt1x7pT1xKH8KfDCOOp2jsfOh
ZpvOMtoiuHH0jTUD47sCFezVXHCgwaK0aczLhjziVvI2D4SICeYVD6yPWyqnneqBA0nrA+iKTMGx
FZ+JGeHlHncJoHwok58rZB+f4s6+X4m4OfKl27jPOd+ijTuUvtHPyozdl8atiiJj7vdbzGXENADy
aNJLUyuU6egqIeVRPbwYqE6NgvNH8VnpVHf0LJpK2BMtyiWvKAM0wU7ir6TrXuFLz981xPbACZVp
9TF6lxWRUS2gBsCT6hb0aOFSXLez0emGIEZ0zesmI4FpV+SVFHA7G1DviBi7sGGGFZYGu3CPvBOo
FvrTBhRMbThA1+dBE0hKEeqfEyVdwkyN+Q7OSNX+VmIk3VrOIstR9qZXZX6hh5HBTRDigYYoIyKc
vftbjUijIocKgekuAHWtSWYTRRQ0yokDCe9O/hckVlVP7m+DRlarZso8orWjQI//IyJ4BZETJnZt
kdCdyobFC9VkNxFtvR0/o4XEO54Ukqrdf18kc54nbTRmn7GQomWOTPTu6FRhcbToey299JZhOoTk
y0FvaRvB0uA1Uo76qMevwkKwvW2fAoHP9otjkYLkfOv85MbJgsaIHzFS2NDIrMV1QWxsBzMQ6pgZ
QpkIWaFb3V2hsvsTvQQXxAZRPx41nLhaBZxAVWSBFRPBnNL62vfv/Er3eeQKd6YCSCdeOGrkAq1n
RGmiheFPNrTSkKpuGEor3Q2UgB8IKmTV8kB7G3FI2r7xGOQe4cYj0cOyEGpOHaQBuMM3UUL1fD5I
suoWuuvGmVQExTd6svCL5rgo/GBTnDF9j7XJkLmt4EZTFIIqOZl/h7oC9pqO7Dkt3i1duzHHec0E
NJ9paLarIcU8cH2F39OFQb/XY4QLnLloKbPSDSVciT86FfRB74xqb96BQx9OuDeuNLEKsvTrORQr
ntMe7jVPZZTsXMX5hFc8KY46hJRUWA+wnGOoPdF4rkoWGp/mFAAZNZ2H3t0vp/s22I9iemfYxvAe
g0lc6wPm0jW3CpdUbvPmBmRUogXIh4vsq/uHUt6ZgMzq490xT2njz9edJdLg3yq2taNgMQW/ty8B
JWp/BFwRcccT5A0CKv7r3RxldCkvWJM5fkMwWzcklC3AvzYAdQ9jE8JS/XjUKr7mbFqWnfSxSoKs
xLKqBDvYOQ0SFAFqJkNOQ6leXX+lHhhjbatSZWChqzoFCLV/ie0Nqr3X9K5X0O72Lk7chWaYilOA
a+1INaCGH+jPk/dMSKx4W2eZxr5b/B9L1Qw2CRwYpovLNTvVDnIvm7VsRH7NPZx/d97yEK+kSPdZ
MhVRRD1HBYe2UH6xbBK1q0UTRg29Ew9oTDD25Zj+ML4bwqd+ypL1ReLZ6Y0MafKu5IrmxN0VdR74
cJbMYZNTwzdNZn40b/vo0+VECptdNJ9lz4Ll7nasp+EPBVuclRKLrzoa/B9Gp6y80hJJxGCPGyCz
e4ICp0xxifVG8+HLvcm9ya54DBWcW/s4mMTe3cm4/CqICjCcq24Z1mGa9RPlQNxNd3b+ANHAbzsi
RgmJAaPpXVLsuv6+MVPvATnWVBwpgp7SS7PcfUNFerM1nLHl0y+g5iaOWStCh2SXtn0fy5dujogC
BSCWF5Eiy6+/qVfx/ndN4/gMnU+6Cb4Pl7hI+92mF4RfD/7SSutYwqOQDnmI9hnCiBHYUFi4eNnB
kR4LXCMurzk5z8hZD5Ud2cRmR+N90pbsIuzlSldqu187/YFV6mcQY9FllIjdlRlqktcFoGQ3Du9Q
cBGSeTgUrcrn4+Zt1z7hv45XOtU3EEzxdfRgqVw3ZFh3D8wpTmD/JcjMuP8IauKbRU2LMlEbqlTp
dki5bjSE557hf7waTrXZ76+K/4HIIXGiG1ObLT+t8Bs3TSmCKMIB+5mKIXXumpr1TCfnWmSAY6hw
+MQE540tQ60sKkYtWw7kK5NzURs1UFmaNMBlGtob3oYIVmRGgzNZ+klMZlHXz5mxO7BCvh1YPZxp
9U+ngq+oEVLyb0AHh6FFNvNR8ygznrPcM9fFeLntCPRWzx+N95D8Px3mGaz5hsT1cKKyN8cZksyj
R96ACpl59g5vvVZ6t53Jsahti93cCi4UVAXFzTfSTQMGsh8j2DfZ4Y714Xa729LcxFlJRzBHSFYs
e0Kd5BzHASHddvTfehzdLZz81Yw4x/av7sEz8/yKUh5v7ZuEa9dFIA4RCLcSID5X/dUTMX2v0SkA
5Le/p9HEuEO71NsDHO82a02kszuduBqZDq/N/6MEyaKKnRw+wNsTjldxbHO2lKrdmc5nmjvqdQmd
qkcTp/WFXXupCkf7tpAAckVqowU30vUGwb9Shn6tePkDKXokJ3NAchLxL7TM2gWUT3AVzorvvjXu
P4vQeEGaho3n+Sf+vAYXC/YURw3Uxf+B8r8fnWKhjMKfm8vMjoRwUbusFxF0Q4DV6IxyB+1iwRAr
mS1eguNc+r1wIr0CE/UKoYENiZYbJtZLa6JScvw4k3CgZN76qAtoLpS7N6xEtcbxZ2M6JEMLBjPg
VWRq6YxmMvhjptOrcrSKGczuzlpqkM3+du3Ew5NTs3V9uyRINHVKjm3YGJJv0QGLbyuffpKm2ZZT
Cwe3hTwyzFyxBR2qddm2EkCTzcJSD/G3Go9QRtArpiXp+bomY736d9+S2N4+3C1oCpM6v62L4+CE
v94EQpc8ajcawZw8yZpRKn8ncPRHCCmMc0jH9kvVZ1e6Ude62jHRKK2AKxoWZxaaDsh4DJ5/1AUZ
KhfyUYKTe5gH+DSb1Yk862JolifuORCHwog9WGv/HOezRzaFisZYTFIovzHb2PTu8NkbkTImkheh
AMqXsZxt9uc20eZRMgZBvavQQXAEBMTmWMM4/BrpRlRhnR4q9G2+zEBdfIrr39QnTiNM1iQ20uoX
xlNfwaVOe6IQb7tA/GVkFmXs/3SNZivAuIUZs51jB5vNp4zy25PpIBuKJSfCQO+b6EbQLUferq9Z
IXazHhMC+s6xGdc/8n4R1CfwOnNhRyCkz5L2kZWKDgOfib2gwcMZD3tVAKSYuqQG3sM3zKNOEdWz
IGVLr4KPWTK4oDm4FbtlNJ/opC9laWf9yu6wnL3PYFFv3OEr9WhHoFe6/ZXoTYN4ZYMphuUvRqYj
qCW4Uq5vINOWDsODJjp47fHrBVtT3oCHPZb9MoGKye5MuLp0xxnnWDTVOAqxChepVntgs5DF1wbX
At/0vUox7WK3ar0zvhBNH35JMvgdTuEXks5HSG4BZZyWNuMoEVSeocA0hN+kBS0veBcRaFnS/M8k
oeXX1YMu8cv2ehcUf9/ouYmMNngrDFg+eSNIdz8bkTZjNBQPMctX7GP/MM5s6tNjuC8OPqGS7eli
d98Vn9m+ip/8gZwep0ZQ7Ddpn4gL4pgCm2FlIKMXSSbj0rWhhFAJpdiSQNcbxRaQhWlHdjbmUmvb
ZMYv5T1pi8kz7LAyzA3ltgvSakQ2rdVUN5+Zd//rTR+3IN7QSIwK5pr8qhAEtCvwFFvy/BmIHsXd
1zuCx4mPB2DnkBaTAjWavFg26fyCO4hxraU1ORbVqs3jxioiJqpHg9I1CQkuG9gYSppO8J7VM4Ms
DvwNIm4CeIJn0J/ii8nIzhpOl31QlQakPheveomAGD8eWPkFt/82NkpkXHf1SC5NMt3WfC6F327i
qw7p8kqxwawRdq8lqkId3zkp15HZCVAmsfc9x5LXQ0/XVZTmmPY2V9qskU94cabOTlUF8jBsPJvv
K1y2+pPqX/B0eZ/U+M13jusuyzr3FhpgfDYXAS6ubCfxqbhpz49WfLoXKj4LgbfYLbpiOsQLm8Vo
qCM5QepHhUJpX90NeDAFqGOOBFbv31Wd5+rsUeqVMsksB9+g0w==

`pragma protect end_protected

endmodule