----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Sun Jan 26 17:25:48 2020
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 19;
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 16;
end coreparameters;
