
-- This is an automatically generated file

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

package coreparameters IS
  constant ARCHITECT : integer := 1;
  constant MODE      : integer := 2;
  constant DP_OPTION : integer := 0;
  constant DP_WIDTH  : integer := 16;
  constant IN_BITS   : integer := 10;
  constant OUT_BITS  : integer := 10;
  constant ROUND     : integer := 1;
  constant COARSE    : integer := 0;
  constant ITERATIONS: integer := 48;
end coreparameters;
