case g_data_samples_exp is
	when 2 =>
		out_cos := (
			to_signed(255, 9), to_signed(0, 9), 
		);
	when 3 =>
		out_cos := (
			to_signed(255, 9), to_signed(180, 9), to_signed(0, 9), to_signed(-180, 9), 
		);
	when 4 =>
		out_cos := (
			to_signed(255, 9), to_signed(236, 9), to_signed(180, 9), to_signed(98, 9), to_signed(0, 9), to_signed(-98, 9), to_signed(-180, 9), to_signed(-236, 9), 
		);
	when 5 =>
		out_cos := (
			to_signed(255, 9), to_signed(250, 9), to_signed(236, 9), to_signed(212, 9), to_signed(180, 9), to_signed(142, 9), to_signed(98, 9), to_signed(50, 9), to_signed(0, 9), to_signed(-50, 9), to_signed(-98, 9), to_signed(-142, 9), to_signed(-180, 9), to_signed(-212, 9), to_signed(-236, 9), to_signed(-250, 9), 
		);
	when 6 =>
		out_cos := (
			to_signed(255, 9), to_signed(254, 9), to_signed(250, 9), to_signed(244, 9), to_signed(236, 9), to_signed(225, 9), to_signed(212, 9), to_signed(197, 9), to_signed(180, 9), to_signed(162, 9), to_signed(142, 9), to_signed(120, 9), to_signed(98, 9), to_signed(74, 9), to_signed(50, 9), to_signed(25, 9), to_signed(0, 9), to_signed(-25, 9), to_signed(-50, 9), to_signed(-74, 9), to_signed(-98, 9), to_signed(-120, 9), to_signed(-142, 9), to_signed(-162, 9), to_signed(-180, 9), to_signed(-197, 9), to_signed(-212, 9), to_signed(-225, 9), to_signed(-236, 9), to_signed(-244, 9), to_signed(-250, 9), to_signed(-254, 9), 
		);
	when 7 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(252, 9), to_signed(250, 9), to_signed(247, 9), to_signed(244, 9), to_signed(240, 9), to_signed(236, 9), to_signed(231, 9), to_signed(225, 9), to_signed(219, 9), to_signed(212, 9), to_signed(205, 9), to_signed(197, 9), to_signed(189, 9), to_signed(180, 9), to_signed(171, 9), to_signed(162, 9), to_signed(152, 9), to_signed(142, 9), to_signed(131, 9), to_signed(120, 9), to_signed(109, 9), to_signed(98, 9), to_signed(86, 9), to_signed(74, 9), to_signed(62, 9), to_signed(50, 9), to_signed(37, 9), to_signed(25, 9), to_signed(13, 9), to_signed(0, 9), to_signed(-13, 9), to_signed(-25, 9), to_signed(-37, 9), to_signed(-50, 9), to_signed(-62, 9), to_signed(-74, 9), to_signed(-86, 9), to_signed(-98, 9), to_signed(-109, 9), to_signed(-120, 9), to_signed(-131, 9), to_signed(-142, 9), to_signed(-152, 9), to_signed(-162, 9), to_signed(-171, 9), to_signed(-180, 9), to_signed(-189, 9), to_signed(-197, 9), to_signed(-205, 9), to_signed(-212, 9), to_signed(-219, 9), to_signed(-225, 9), to_signed(-231, 9), to_signed(-236, 9), to_signed(-240, 9), to_signed(-244, 9), to_signed(-247, 9), to_signed(-250, 9), to_signed(-252, 9), to_signed(-254, 9), to_signed(-255, 9), 
		);
	when 8 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(252, 9), to_signed(251, 9), to_signed(250, 9), to_signed(249, 9), to_signed(247, 9), to_signed(246, 9), to_signed(244, 9), to_signed(242, 9), to_signed(240, 9), to_signed(238, 9), to_signed(236, 9), to_signed(233, 9), to_signed(231, 9), to_signed(228, 9), to_signed(225, 9), to_signed(222, 9), to_signed(219, 9), to_signed(215, 9), to_signed(212, 9), to_signed(208, 9), to_signed(205, 9), to_signed(201, 9), to_signed(197, 9), to_signed(193, 9), to_signed(189, 9), to_signed(185, 9), to_signed(180, 9), to_signed(176, 9), to_signed(171, 9), to_signed(167, 9), to_signed(162, 9), to_signed(157, 9), to_signed(152, 9), to_signed(147, 9), to_signed(142, 9), to_signed(136, 9), to_signed(131, 9), to_signed(126, 9), to_signed(120, 9), to_signed(115, 9), to_signed(109, 9), to_signed(103, 9), to_signed(98, 9), to_signed(92, 9), to_signed(86, 9), to_signed(80, 9), to_signed(74, 9), to_signed(68, 9), to_signed(62, 9), to_signed(56, 9), to_signed(50, 9), to_signed(44, 9), to_signed(37, 9), to_signed(31, 9), to_signed(25, 9), to_signed(19, 9), to_signed(13, 9), to_signed(6, 9), to_signed(0, 9), to_signed(-6, 9), to_signed(-13, 9), to_signed(-19, 9), to_signed(-25, 9), to_signed(-31, 9), to_signed(-37, 9), to_signed(-44, 9), to_signed(-50, 9), to_signed(-56, 9), to_signed(-62, 9), to_signed(-68, 9), to_signed(-74, 9), to_signed(-80, 9), to_signed(-86, 9), to_signed(-92, 9), to_signed(-98, 9), to_signed(-103, 9), to_signed(-109, 9), to_signed(-115, 9), to_signed(-120, 9), to_signed(-126, 9), to_signed(-131, 9), to_signed(-136, 9), to_signed(-142, 9), to_signed(-147, 9), to_signed(-152, 9), to_signed(-157, 9), to_signed(-162, 9), to_signed(-167, 9), to_signed(-171, 9), to_signed(-176, 9), to_signed(-180, 9), to_signed(-185, 9), to_signed(-189, 9), to_signed(-193, 9), to_signed(-197, 9), to_signed(-201, 9), to_signed(-205, 9), to_signed(-208, 9), to_signed(-212, 9), to_signed(-215, 9), to_signed(-219, 9), to_signed(-222, 9), to_signed(-225, 9), to_signed(-228, 9), to_signed(-231, 9), to_signed(-233, 9), to_signed(-236, 9), to_signed(-238, 9), to_signed(-240, 9), to_signed(-242, 9), to_signed(-244, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 9 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(245, 9), to_signed(244, 9), to_signed(243, 9), to_signed(242, 9), to_signed(241, 9), to_signed(240, 9), to_signed(239, 9), to_signed(238, 9), to_signed(237, 9), to_signed(236, 9), to_signed(234, 9), to_signed(233, 9), to_signed(232, 9), to_signed(231, 9), to_signed(229, 9), to_signed(228, 9), to_signed(226, 9), to_signed(225, 9), to_signed(223, 9), to_signed(222, 9), to_signed(220, 9), to_signed(219, 9), to_signed(217, 9), to_signed(215, 9), to_signed(214, 9), to_signed(212, 9), to_signed(210, 9), to_signed(208, 9), to_signed(207, 9), to_signed(205, 9), to_signed(203, 9), to_signed(201, 9), to_signed(199, 9), to_signed(197, 9), to_signed(195, 9), to_signed(193, 9), to_signed(191, 9), to_signed(189, 9), to_signed(187, 9), to_signed(185, 9), to_signed(183, 9), to_signed(180, 9), to_signed(178, 9), to_signed(176, 9), to_signed(174, 9), to_signed(171, 9), to_signed(169, 9), to_signed(167, 9), to_signed(164, 9), to_signed(162, 9), to_signed(159, 9), to_signed(157, 9), to_signed(154, 9), to_signed(152, 9), to_signed(149, 9), to_signed(147, 9), to_signed(144, 9), to_signed(142, 9), to_signed(139, 9), to_signed(136, 9), to_signed(134, 9), to_signed(131, 9), to_signed(128, 9), to_signed(126, 9), to_signed(123, 9), to_signed(120, 9), to_signed(117, 9), to_signed(115, 9), to_signed(112, 9), to_signed(109, 9), to_signed(106, 9), to_signed(103, 9), to_signed(100, 9), to_signed(98, 9), to_signed(95, 9), to_signed(92, 9), to_signed(89, 9), to_signed(86, 9), to_signed(83, 9), to_signed(80, 9), to_signed(77, 9), to_signed(74, 9), to_signed(71, 9), to_signed(68, 9), to_signed(65, 9), to_signed(62, 9), to_signed(59, 9), to_signed(56, 9), to_signed(53, 9), to_signed(50, 9), to_signed(47, 9), to_signed(44, 9), to_signed(41, 9), to_signed(37, 9), to_signed(34, 9), to_signed(31, 9), to_signed(28, 9), to_signed(25, 9), to_signed(22, 9), to_signed(19, 9), to_signed(16, 9), to_signed(13, 9), to_signed(9, 9), to_signed(6, 9), to_signed(3, 9), to_signed(0, 9), to_signed(-3, 9), to_signed(-6, 9), to_signed(-9, 9), to_signed(-13, 9), to_signed(-16, 9), to_signed(-19, 9), to_signed(-22, 9), to_signed(-25, 9), to_signed(-28, 9), to_signed(-31, 9), to_signed(-34, 9), to_signed(-37, 9), to_signed(-41, 9), to_signed(-44, 9), to_signed(-47, 9), to_signed(-50, 9), to_signed(-53, 9), to_signed(-56, 9), to_signed(-59, 9), to_signed(-62, 9), to_signed(-65, 9), to_signed(-68, 9), to_signed(-71, 9), to_signed(-74, 9), to_signed(-77, 9), to_signed(-80, 9), to_signed(-83, 9), to_signed(-86, 9), to_signed(-89, 9), to_signed(-92, 9), to_signed(-95, 9), to_signed(-98, 9), to_signed(-100, 9), to_signed(-103, 9), to_signed(-106, 9), to_signed(-109, 9), to_signed(-112, 9), to_signed(-115, 9), to_signed(-117, 9), to_signed(-120, 9), to_signed(-123, 9), to_signed(-126, 9), to_signed(-128, 9), to_signed(-131, 9), to_signed(-134, 9), to_signed(-136, 9), to_signed(-139, 9), to_signed(-142, 9), to_signed(-144, 9), to_signed(-147, 9), to_signed(-149, 9), to_signed(-152, 9), to_signed(-154, 9), to_signed(-157, 9), to_signed(-159, 9), to_signed(-162, 9), to_signed(-164, 9), to_signed(-167, 9), to_signed(-169, 9), to_signed(-171, 9), to_signed(-174, 9), to_signed(-176, 9), to_signed(-178, 9), to_signed(-180, 9), to_signed(-183, 9), to_signed(-185, 9), to_signed(-187, 9), to_signed(-189, 9), to_signed(-191, 9), to_signed(-193, 9), to_signed(-195, 9), to_signed(-197, 9), to_signed(-199, 9), to_signed(-201, 9), to_signed(-203, 9), to_signed(-205, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-210, 9), to_signed(-212, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-217, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 10 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(218, 9), to_signed(217, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(213, 9), to_signed(212, 9), to_signed(211, 9), to_signed(210, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(206, 9), to_signed(205, 9), to_signed(204, 9), to_signed(203, 9), to_signed(202, 9), to_signed(201, 9), to_signed(200, 9), to_signed(199, 9), to_signed(198, 9), to_signed(197, 9), to_signed(196, 9), to_signed(195, 9), to_signed(194, 9), to_signed(193, 9), to_signed(192, 9), to_signed(191, 9), to_signed(190, 9), to_signed(189, 9), to_signed(188, 9), to_signed(187, 9), to_signed(186, 9), to_signed(185, 9), to_signed(184, 9), to_signed(183, 9), to_signed(181, 9), to_signed(180, 9), to_signed(179, 9), to_signed(178, 9), to_signed(177, 9), to_signed(176, 9), to_signed(175, 9), to_signed(174, 9), to_signed(172, 9), to_signed(171, 9), to_signed(170, 9), to_signed(169, 9), to_signed(168, 9), to_signed(167, 9), to_signed(165, 9), to_signed(164, 9), to_signed(163, 9), to_signed(162, 9), to_signed(161, 9), to_signed(159, 9), to_signed(158, 9), to_signed(157, 9), to_signed(156, 9), to_signed(154, 9), to_signed(153, 9), to_signed(152, 9), to_signed(151, 9), to_signed(149, 9), to_signed(148, 9), to_signed(147, 9), to_signed(146, 9), to_signed(144, 9), to_signed(143, 9), to_signed(142, 9), to_signed(140, 9), to_signed(139, 9), to_signed(138, 9), to_signed(136, 9), to_signed(135, 9), to_signed(134, 9), to_signed(132, 9), to_signed(131, 9), to_signed(130, 9), to_signed(128, 9), to_signed(127, 9), to_signed(126, 9), to_signed(124, 9), to_signed(123, 9), to_signed(122, 9), to_signed(120, 9), to_signed(119, 9), to_signed(117, 9), to_signed(116, 9), to_signed(115, 9), to_signed(113, 9), to_signed(112, 9), to_signed(110, 9), to_signed(109, 9), to_signed(108, 9), to_signed(106, 9), to_signed(105, 9), to_signed(103, 9), to_signed(102, 9), to_signed(100, 9), to_signed(99, 9), to_signed(98, 9), to_signed(96, 9), to_signed(95, 9), to_signed(93, 9), to_signed(92, 9), to_signed(90, 9), to_signed(89, 9), to_signed(87, 9), to_signed(86, 9), to_signed(84, 9), to_signed(83, 9), to_signed(81, 9), to_signed(80, 9), to_signed(79, 9), to_signed(77, 9), to_signed(76, 9), to_signed(74, 9), to_signed(73, 9), to_signed(71, 9), to_signed(70, 9), to_signed(68, 9), to_signed(67, 9), to_signed(65, 9), to_signed(63, 9), to_signed(62, 9), to_signed(60, 9), to_signed(59, 9), to_signed(57, 9), to_signed(56, 9), to_signed(54, 9), to_signed(53, 9), to_signed(51, 9), to_signed(50, 9), to_signed(48, 9), to_signed(47, 9), to_signed(45, 9), to_signed(44, 9), to_signed(42, 9), to_signed(41, 9), to_signed(39, 9), to_signed(37, 9), to_signed(36, 9), to_signed(34, 9), to_signed(33, 9), to_signed(31, 9), to_signed(30, 9), to_signed(28, 9), to_signed(27, 9), to_signed(25, 9), to_signed(23, 9), to_signed(22, 9), to_signed(20, 9), to_signed(19, 9), to_signed(17, 9), to_signed(16, 9), to_signed(14, 9), to_signed(13, 9), to_signed(11, 9), to_signed(9, 9), to_signed(8, 9), to_signed(6, 9), to_signed(5, 9), to_signed(3, 9), to_signed(2, 9), to_signed(0, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-11, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-25, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-39, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-65, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 11 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(65, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(49, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(39, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(32, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(25, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(18, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(11, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(7, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 12 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(119, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(112, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(106, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(101, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(97, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(92, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(89, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(85, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(82, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(78, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(75, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(72, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(69, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(66, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(64, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(61, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(58, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(56, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(53, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(50, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(48, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(45, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(43, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(40, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(38, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(36, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(33, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(31, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(29, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(26, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(24, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(22, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(19, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(17, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(15, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(12, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(10, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(8, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(6, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(3, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(1, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 13 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 14 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 15 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when 16 =>
		out_cos := (
			to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(255, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(254, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(253, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(252, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(251, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(250, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(249, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(248, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(247, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(246, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(245, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(244, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(243, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(242, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(241, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(240, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(239, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(238, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(237, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(236, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(235, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(234, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(233, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(232, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(231, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(230, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(229, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(228, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(227, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(226, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(225, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(224, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(223, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(222, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(221, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(220, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(219, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(218, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(217, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(216, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(215, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(214, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(213, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(212, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(211, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(210, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(209, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(208, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(207, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(206, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(205, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(204, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(203, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(202, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(201, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(200, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(199, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(198, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(197, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(196, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(195, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(194, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(193, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(192, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(191, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(190, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(189, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(188, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(187, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(186, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(185, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(184, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(183, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(182, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(181, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(180, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(179, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(178, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(177, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(176, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(175, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(174, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(173, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(172, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(171, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(170, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(169, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(168, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(167, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(166, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(165, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(164, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(163, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(162, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(161, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(160, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(159, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(158, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(157, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(156, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(155, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(154, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(153, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(152, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(151, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(150, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(149, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(148, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(147, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(146, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(145, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(144, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(143, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(142, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(141, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(140, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(139, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(138, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(137, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(136, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(135, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(134, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(133, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(132, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(131, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(130, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(129, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(128, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(127, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(126, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(125, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(124, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(123, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(122, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(121, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(120, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(119, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(118, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(117, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(116, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(115, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(114, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(113, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(112, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(111, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(110, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(109, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(108, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(107, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(106, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(105, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(104, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(103, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(102, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(101, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(100, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(99, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(98, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(97, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(96, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(95, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(94, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(93, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(92, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(91, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(90, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(89, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(88, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(87, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(86, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(85, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(84, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(83, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(82, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(81, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(80, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(79, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(78, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(77, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(76, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(75, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(74, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(73, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(72, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(71, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(70, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(69, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(68, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(67, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(66, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(65, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(64, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(63, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(62, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(61, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(60, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(59, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(58, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(57, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(56, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(55, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(54, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(53, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(52, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(51, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(50, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(49, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(48, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(47, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(46, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(45, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(44, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(43, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(42, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(41, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(40, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(39, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(38, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(37, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(36, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(35, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(34, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(33, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(32, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(31, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(30, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(29, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(28, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(27, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(26, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(25, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(24, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(23, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(22, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(21, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(20, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(19, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(18, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(17, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(16, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(15, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(14, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(13, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(12, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(11, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(10, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(9, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(8, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(7, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(6, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(5, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(4, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(3, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(2, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(1, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(0, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-1, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-2, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-3, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-4, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-5, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-6, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-7, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-8, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-9, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-10, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-11, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-12, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-13, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-14, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-15, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-16, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-17, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-18, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-19, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-20, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-21, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-22, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-23, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-24, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-25, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-26, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-27, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-28, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-29, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-30, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-31, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-32, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-33, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-34, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-35, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-36, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-37, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-38, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-39, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-40, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-41, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-42, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-43, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-44, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-45, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-46, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-47, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-48, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-49, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-50, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-51, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-52, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-53, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-54, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-55, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-56, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-57, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-58, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-59, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-60, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-61, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-62, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-63, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-64, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-65, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-66, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-67, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-68, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-69, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-70, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-71, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-72, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-73, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-74, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-75, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-76, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-77, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-78, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-79, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-80, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-81, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-82, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-83, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-84, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-85, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-86, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-87, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-88, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-89, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-90, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-91, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-92, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-93, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-94, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-95, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-96, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-97, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-98, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-99, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-100, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-101, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-102, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-103, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-104, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-105, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-106, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-107, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-108, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-109, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-110, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-111, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-112, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-113, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-114, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-115, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-116, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-117, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-118, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-119, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-120, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-121, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-122, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-123, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-124, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-125, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-126, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-127, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-128, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-129, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-130, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-131, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-132, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-133, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-134, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-135, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-136, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-137, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-138, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-139, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-140, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-141, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-142, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-143, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-144, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-145, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-146, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-147, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-148, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-149, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-150, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-151, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-152, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-153, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-154, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-155, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-156, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-157, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-158, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-159, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-160, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-161, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-162, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-163, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-164, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-165, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-166, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-167, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-168, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-169, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-170, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-171, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-172, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-173, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-174, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-175, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-176, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-177, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-178, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-179, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-180, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-181, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-182, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-183, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-184, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-185, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-186, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-187, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-188, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-189, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-190, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-191, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-192, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-193, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-194, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-195, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-196, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-197, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-198, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-199, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-200, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-201, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-202, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-203, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-204, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-205, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-206, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-207, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-208, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-209, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-210, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-211, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-212, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-213, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-214, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-215, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-216, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-217, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-218, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-219, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-220, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-221, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-222, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-223, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-224, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-225, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-226, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-227, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-228, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-229, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-230, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-231, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-232, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-233, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-234, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-235, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-236, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-237, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-238, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-239, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-240, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-241, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-242, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-243, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-244, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-245, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-246, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-247, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-248, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-249, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-250, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-251, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-252, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-253, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-254, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), to_signed(-255, 9), 
		);
	when others =>
		out_cos := (others => "011111111");
end case;